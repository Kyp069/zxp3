
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"1c",x"00",x"00",x"36"),
     1 => (x"41",x"41",x"63",x"3e"),
     2 => (x"7f",x"00",x"00",x"41"),
     3 => (x"3e",x"63",x"41",x"7f"),
     4 => (x"7f",x"00",x"00",x"1c"),
     5 => (x"41",x"49",x"49",x"7f"),
     6 => (x"7f",x"00",x"00",x"41"),
     7 => (x"01",x"09",x"09",x"7f"),
     8 => (x"3e",x"00",x"00",x"01"),
     9 => (x"7b",x"49",x"41",x"7f"),
    10 => (x"7f",x"00",x"00",x"7a"),
    11 => (x"7f",x"08",x"08",x"7f"),
    12 => (x"00",x"00",x"00",x"7f"),
    13 => (x"41",x"7f",x"7f",x"41"),
    14 => (x"20",x"00",x"00",x"00"),
    15 => (x"7f",x"40",x"40",x"60"),
    16 => (x"7f",x"7f",x"00",x"3f"),
    17 => (x"63",x"36",x"1c",x"08"),
    18 => (x"7f",x"00",x"00",x"41"),
    19 => (x"40",x"40",x"40",x"7f"),
    20 => (x"7f",x"7f",x"00",x"40"),
    21 => (x"7f",x"06",x"0c",x"06"),
    22 => (x"7f",x"7f",x"00",x"7f"),
    23 => (x"7f",x"18",x"0c",x"06"),
    24 => (x"3e",x"00",x"00",x"7f"),
    25 => (x"7f",x"41",x"41",x"7f"),
    26 => (x"7f",x"00",x"00",x"3e"),
    27 => (x"0f",x"09",x"09",x"7f"),
    28 => (x"7f",x"3e",x"00",x"06"),
    29 => (x"7e",x"7f",x"61",x"41"),
    30 => (x"7f",x"00",x"00",x"40"),
    31 => (x"7f",x"19",x"09",x"7f"),
    32 => (x"26",x"00",x"00",x"66"),
    33 => (x"7b",x"59",x"4d",x"6f"),
    34 => (x"01",x"00",x"00",x"32"),
    35 => (x"01",x"7f",x"7f",x"01"),
    36 => (x"3f",x"00",x"00",x"01"),
    37 => (x"7f",x"40",x"40",x"7f"),
    38 => (x"0f",x"00",x"00",x"3f"),
    39 => (x"3f",x"70",x"70",x"3f"),
    40 => (x"7f",x"7f",x"00",x"0f"),
    41 => (x"7f",x"30",x"18",x"30"),
    42 => (x"63",x"41",x"00",x"7f"),
    43 => (x"36",x"1c",x"1c",x"36"),
    44 => (x"03",x"01",x"41",x"63"),
    45 => (x"06",x"7c",x"7c",x"06"),
    46 => (x"71",x"61",x"01",x"03"),
    47 => (x"43",x"47",x"4d",x"59"),
    48 => (x"00",x"00",x"00",x"41"),
    49 => (x"41",x"41",x"7f",x"7f"),
    50 => (x"03",x"01",x"00",x"00"),
    51 => (x"30",x"18",x"0c",x"06"),
    52 => (x"00",x"00",x"40",x"60"),
    53 => (x"7f",x"7f",x"41",x"41"),
    54 => (x"0c",x"08",x"00",x"00"),
    55 => (x"0c",x"06",x"03",x"06"),
    56 => (x"80",x"80",x"00",x"08"),
    57 => (x"80",x"80",x"80",x"80"),
    58 => (x"00",x"00",x"00",x"80"),
    59 => (x"04",x"07",x"03",x"00"),
    60 => (x"20",x"00",x"00",x"00"),
    61 => (x"7c",x"54",x"54",x"74"),
    62 => (x"7f",x"00",x"00",x"78"),
    63 => (x"7c",x"44",x"44",x"7f"),
    64 => (x"38",x"00",x"00",x"38"),
    65 => (x"44",x"44",x"44",x"7c"),
    66 => (x"38",x"00",x"00",x"00"),
    67 => (x"7f",x"44",x"44",x"7c"),
    68 => (x"38",x"00",x"00",x"7f"),
    69 => (x"5c",x"54",x"54",x"7c"),
    70 => (x"04",x"00",x"00",x"18"),
    71 => (x"05",x"05",x"7f",x"7e"),
    72 => (x"18",x"00",x"00",x"00"),
    73 => (x"fc",x"a4",x"a4",x"bc"),
    74 => (x"7f",x"00",x"00",x"7c"),
    75 => (x"7c",x"04",x"04",x"7f"),
    76 => (x"00",x"00",x"00",x"78"),
    77 => (x"40",x"7d",x"3d",x"00"),
    78 => (x"80",x"00",x"00",x"00"),
    79 => (x"7d",x"fd",x"80",x"80"),
    80 => (x"7f",x"00",x"00",x"00"),
    81 => (x"6c",x"38",x"10",x"7f"),
    82 => (x"00",x"00",x"00",x"44"),
    83 => (x"40",x"7f",x"3f",x"00"),
    84 => (x"7c",x"7c",x"00",x"00"),
    85 => (x"7c",x"0c",x"18",x"0c"),
    86 => (x"7c",x"00",x"00",x"78"),
    87 => (x"7c",x"04",x"04",x"7c"),
    88 => (x"38",x"00",x"00",x"78"),
    89 => (x"7c",x"44",x"44",x"7c"),
    90 => (x"fc",x"00",x"00",x"38"),
    91 => (x"3c",x"24",x"24",x"fc"),
    92 => (x"18",x"00",x"00",x"18"),
    93 => (x"fc",x"24",x"24",x"3c"),
    94 => (x"7c",x"00",x"00",x"fc"),
    95 => (x"0c",x"04",x"04",x"7c"),
    96 => (x"48",x"00",x"00",x"08"),
    97 => (x"74",x"54",x"54",x"5c"),
    98 => (x"04",x"00",x"00",x"20"),
    99 => (x"44",x"44",x"7f",x"3f"),
   100 => (x"3c",x"00",x"00",x"00"),
   101 => (x"7c",x"40",x"40",x"7c"),
   102 => (x"1c",x"00",x"00",x"7c"),
   103 => (x"3c",x"60",x"60",x"3c"),
   104 => (x"7c",x"3c",x"00",x"1c"),
   105 => (x"7c",x"60",x"30",x"60"),
   106 => (x"6c",x"44",x"00",x"3c"),
   107 => (x"6c",x"38",x"10",x"38"),
   108 => (x"1c",x"00",x"00",x"44"),
   109 => (x"3c",x"60",x"e0",x"bc"),
   110 => (x"44",x"00",x"00",x"1c"),
   111 => (x"4c",x"5c",x"74",x"64"),
   112 => (x"08",x"00",x"00",x"44"),
   113 => (x"41",x"77",x"3e",x"08"),
   114 => (x"00",x"00",x"00",x"41"),
   115 => (x"00",x"7f",x"7f",x"00"),
   116 => (x"41",x"00",x"00",x"00"),
   117 => (x"08",x"3e",x"77",x"41"),
   118 => (x"01",x"02",x"00",x"08"),
   119 => (x"02",x"02",x"03",x"01"),
   120 => (x"7f",x"7f",x"00",x"01"),
   121 => (x"7f",x"7f",x"7f",x"7f"),
   122 => (x"08",x"08",x"00",x"7f"),
   123 => (x"3e",x"3e",x"1c",x"1c"),
   124 => (x"7f",x"7f",x"7f",x"7f"),
   125 => (x"1c",x"1c",x"3e",x"3e"),
   126 => (x"10",x"00",x"08",x"08"),
   127 => (x"18",x"7c",x"7c",x"18"),
   128 => (x"10",x"00",x"00",x"10"),
   129 => (x"30",x"7c",x"7c",x"30"),
   130 => (x"30",x"10",x"00",x"10"),
   131 => (x"1e",x"78",x"60",x"60"),
   132 => (x"66",x"42",x"00",x"06"),
   133 => (x"66",x"3c",x"18",x"3c"),
   134 => (x"38",x"78",x"00",x"42"),
   135 => (x"6c",x"c6",x"c2",x"6a"),
   136 => (x"00",x"60",x"00",x"38"),
   137 => (x"00",x"00",x"60",x"00"),
   138 => (x"5e",x"0e",x"00",x"60"),
   139 => (x"0e",x"5d",x"5c",x"5b"),
   140 => (x"c2",x"4c",x"71",x"1e"),
   141 => (x"4d",x"bf",x"d9",x"f6"),
   142 => (x"1e",x"c0",x"4b",x"c0"),
   143 => (x"c7",x"02",x"ab",x"74"),
   144 => (x"48",x"a6",x"c4",x"87"),
   145 => (x"87",x"c5",x"78",x"c0"),
   146 => (x"c1",x"48",x"a6",x"c4"),
   147 => (x"1e",x"66",x"c4",x"78"),
   148 => (x"df",x"ee",x"49",x"73"),
   149 => (x"c0",x"86",x"c8",x"87"),
   150 => (x"ef",x"ef",x"49",x"e0"),
   151 => (x"4a",x"a5",x"c4",x"87"),
   152 => (x"f0",x"f0",x"49",x"6a"),
   153 => (x"87",x"c6",x"f1",x"87"),
   154 => (x"83",x"c1",x"85",x"cb"),
   155 => (x"04",x"ab",x"b7",x"c8"),
   156 => (x"26",x"87",x"c7",x"ff"),
   157 => (x"4c",x"26",x"4d",x"26"),
   158 => (x"4f",x"26",x"4b",x"26"),
   159 => (x"c2",x"4a",x"71",x"1e"),
   160 => (x"c2",x"5a",x"dd",x"f6"),
   161 => (x"c7",x"48",x"dd",x"f6"),
   162 => (x"dd",x"fe",x"49",x"78"),
   163 => (x"1e",x"4f",x"26",x"87"),
   164 => (x"4a",x"71",x"1e",x"73"),
   165 => (x"03",x"aa",x"b7",x"c0"),
   166 => (x"d7",x"c2",x"87",x"d3"),
   167 => (x"c4",x"05",x"bf",x"e0"),
   168 => (x"c2",x"4b",x"c1",x"87"),
   169 => (x"c2",x"4b",x"c0",x"87"),
   170 => (x"c4",x"5b",x"e4",x"d7"),
   171 => (x"e4",x"d7",x"c2",x"87"),
   172 => (x"e0",x"d7",x"c2",x"5a"),
   173 => (x"9a",x"c1",x"4a",x"bf"),
   174 => (x"49",x"a2",x"c0",x"c1"),
   175 => (x"fc",x"87",x"e8",x"ec"),
   176 => (x"e0",x"d7",x"c2",x"48"),
   177 => (x"ef",x"fe",x"78",x"bf"),
   178 => (x"4a",x"71",x"1e",x"87"),
   179 => (x"72",x"1e",x"66",x"c4"),
   180 => (x"87",x"ee",x"e9",x"49"),
   181 => (x"1e",x"4f",x"26",x"26"),
   182 => (x"bf",x"e0",x"d7",x"c2"),
   183 => (x"87",x"f3",x"e5",x"49"),
   184 => (x"48",x"d1",x"f6",x"c2"),
   185 => (x"c2",x"78",x"bf",x"e8"),
   186 => (x"ec",x"48",x"cd",x"f6"),
   187 => (x"f6",x"c2",x"78",x"bf"),
   188 => (x"49",x"4a",x"bf",x"d1"),
   189 => (x"c8",x"99",x"ff",x"c3"),
   190 => (x"48",x"72",x"2a",x"b7"),
   191 => (x"f6",x"c2",x"b0",x"71"),
   192 => (x"4f",x"26",x"58",x"d9"),
   193 => (x"5c",x"5b",x"5e",x"0e"),
   194 => (x"4b",x"71",x"0e",x"5d"),
   195 => (x"c2",x"87",x"c8",x"ff"),
   196 => (x"c0",x"48",x"cc",x"f6"),
   197 => (x"e5",x"49",x"73",x"50"),
   198 => (x"49",x"70",x"87",x"d9"),
   199 => (x"cb",x"9c",x"c2",x"4c"),
   200 => (x"c3",x"cb",x"49",x"ee"),
   201 => (x"4d",x"49",x"70",x"87"),
   202 => (x"97",x"cc",x"f6",x"c2"),
   203 => (x"e2",x"c1",x"05",x"bf"),
   204 => (x"49",x"66",x"d0",x"87"),
   205 => (x"bf",x"d5",x"f6",x"c2"),
   206 => (x"87",x"d6",x"05",x"99"),
   207 => (x"c2",x"49",x"66",x"d4"),
   208 => (x"99",x"bf",x"cd",x"f6"),
   209 => (x"73",x"87",x"cb",x"05"),
   210 => (x"87",x"e7",x"e4",x"49"),
   211 => (x"c1",x"02",x"98",x"70"),
   212 => (x"4c",x"c1",x"87",x"c1"),
   213 => (x"75",x"87",x"c0",x"fe"),
   214 => (x"87",x"d8",x"ca",x"49"),
   215 => (x"c6",x"02",x"98",x"70"),
   216 => (x"cc",x"f6",x"c2",x"87"),
   217 => (x"c2",x"50",x"c1",x"48"),
   218 => (x"bf",x"97",x"cc",x"f6"),
   219 => (x"87",x"e3",x"c0",x"05"),
   220 => (x"bf",x"d5",x"f6",x"c2"),
   221 => (x"99",x"66",x"d0",x"49"),
   222 => (x"87",x"d6",x"ff",x"05"),
   223 => (x"bf",x"cd",x"f6",x"c2"),
   224 => (x"99",x"66",x"d4",x"49"),
   225 => (x"87",x"ca",x"ff",x"05"),
   226 => (x"e6",x"e3",x"49",x"73"),
   227 => (x"05",x"98",x"70",x"87"),
   228 => (x"74",x"87",x"ff",x"fe"),
   229 => (x"87",x"dc",x"fb",x"48"),
   230 => (x"5c",x"5b",x"5e",x"0e"),
   231 => (x"86",x"f4",x"0e",x"5d"),
   232 => (x"ec",x"4c",x"4d",x"c0"),
   233 => (x"a6",x"c4",x"7e",x"bf"),
   234 => (x"d9",x"f6",x"c2",x"48"),
   235 => (x"1e",x"c1",x"78",x"bf"),
   236 => (x"49",x"c7",x"1e",x"c0"),
   237 => (x"c8",x"87",x"cd",x"fd"),
   238 => (x"02",x"98",x"70",x"86"),
   239 => (x"49",x"ff",x"87",x"cd"),
   240 => (x"c1",x"87",x"cc",x"fb"),
   241 => (x"ea",x"e2",x"49",x"da"),
   242 => (x"c2",x"4d",x"c1",x"87"),
   243 => (x"bf",x"97",x"cc",x"f6"),
   244 => (x"cf",x"87",x"c3",x"02"),
   245 => (x"f6",x"c2",x"87",x"fc"),
   246 => (x"c2",x"4b",x"bf",x"d1"),
   247 => (x"05",x"bf",x"e0",x"d7"),
   248 => (x"c3",x"87",x"e9",x"c0"),
   249 => (x"ca",x"e2",x"49",x"fd"),
   250 => (x"49",x"fa",x"c3",x"87"),
   251 => (x"73",x"87",x"c4",x"e2"),
   252 => (x"99",x"ff",x"c3",x"49"),
   253 => (x"49",x"c0",x"1e",x"71"),
   254 => (x"73",x"87",x"ce",x"fb"),
   255 => (x"29",x"b7",x"c8",x"49"),
   256 => (x"49",x"c1",x"1e",x"71"),
   257 => (x"c8",x"87",x"c2",x"fb"),
   258 => (x"87",x"fa",x"c5",x"86"),
   259 => (x"bf",x"d5",x"f6",x"c2"),
   260 => (x"dd",x"02",x"9b",x"4b"),
   261 => (x"dc",x"d7",x"c2",x"87"),
   262 => (x"d7",x"c7",x"49",x"bf"),
   263 => (x"05",x"98",x"70",x"87"),
   264 => (x"4b",x"c0",x"87",x"c4"),
   265 => (x"e0",x"c2",x"87",x"d2"),
   266 => (x"87",x"fc",x"c6",x"49"),
   267 => (x"58",x"e0",x"d7",x"c2"),
   268 => (x"d7",x"c2",x"87",x"c6"),
   269 => (x"78",x"c0",x"48",x"dc"),
   270 => (x"99",x"c2",x"49",x"73"),
   271 => (x"c3",x"87",x"cd",x"05"),
   272 => (x"ee",x"e0",x"49",x"eb"),
   273 => (x"c2",x"49",x"70",x"87"),
   274 => (x"87",x"c2",x"02",x"99"),
   275 => (x"49",x"73",x"4c",x"fb"),
   276 => (x"cd",x"05",x"99",x"c1"),
   277 => (x"49",x"f4",x"c3",x"87"),
   278 => (x"70",x"87",x"d8",x"e0"),
   279 => (x"02",x"99",x"c2",x"49"),
   280 => (x"4c",x"fa",x"87",x"c2"),
   281 => (x"99",x"c8",x"49",x"73"),
   282 => (x"c3",x"87",x"cd",x"05"),
   283 => (x"c2",x"e0",x"49",x"f5"),
   284 => (x"c2",x"49",x"70",x"87"),
   285 => (x"87",x"d4",x"02",x"99"),
   286 => (x"bf",x"dd",x"f6",x"c2"),
   287 => (x"48",x"87",x"c9",x"02"),
   288 => (x"f6",x"c2",x"88",x"c1"),
   289 => (x"87",x"c2",x"58",x"e1"),
   290 => (x"4d",x"c1",x"4c",x"ff"),
   291 => (x"99",x"c4",x"49",x"73"),
   292 => (x"c3",x"87",x"ce",x"05"),
   293 => (x"df",x"ff",x"49",x"f2"),
   294 => (x"49",x"70",x"87",x"d9"),
   295 => (x"db",x"02",x"99",x"c2"),
   296 => (x"dd",x"f6",x"c2",x"87"),
   297 => (x"c7",x"48",x"7e",x"bf"),
   298 => (x"cb",x"03",x"a8",x"b7"),
   299 => (x"c1",x"48",x"6e",x"87"),
   300 => (x"e1",x"f6",x"c2",x"80"),
   301 => (x"87",x"c2",x"c0",x"58"),
   302 => (x"4d",x"c1",x"4c",x"fe"),
   303 => (x"ff",x"49",x"fd",x"c3"),
   304 => (x"70",x"87",x"f0",x"de"),
   305 => (x"02",x"99",x"c2",x"49"),
   306 => (x"f6",x"c2",x"87",x"d5"),
   307 => (x"c0",x"02",x"bf",x"dd"),
   308 => (x"f6",x"c2",x"87",x"c9"),
   309 => (x"78",x"c0",x"48",x"dd"),
   310 => (x"fd",x"87",x"c2",x"c0"),
   311 => (x"c3",x"4d",x"c1",x"4c"),
   312 => (x"de",x"ff",x"49",x"fa"),
   313 => (x"49",x"70",x"87",x"cd"),
   314 => (x"d9",x"02",x"99",x"c2"),
   315 => (x"dd",x"f6",x"c2",x"87"),
   316 => (x"b7",x"c7",x"48",x"bf"),
   317 => (x"c9",x"c0",x"03",x"a8"),
   318 => (x"dd",x"f6",x"c2",x"87"),
   319 => (x"c0",x"78",x"c7",x"48"),
   320 => (x"4c",x"fc",x"87",x"c2"),
   321 => (x"b7",x"c0",x"4d",x"c1"),
   322 => (x"d1",x"c0",x"03",x"ac"),
   323 => (x"4a",x"66",x"c4",x"87"),
   324 => (x"6a",x"82",x"d8",x"c1"),
   325 => (x"87",x"c6",x"c0",x"02"),
   326 => (x"49",x"74",x"4b",x"6a"),
   327 => (x"1e",x"c0",x"0f",x"73"),
   328 => (x"c1",x"1e",x"f0",x"c3"),
   329 => (x"db",x"f7",x"49",x"da"),
   330 => (x"70",x"86",x"c8",x"87"),
   331 => (x"e2",x"c0",x"02",x"98"),
   332 => (x"48",x"a6",x"c8",x"87"),
   333 => (x"bf",x"dd",x"f6",x"c2"),
   334 => (x"49",x"66",x"c8",x"78"),
   335 => (x"66",x"c4",x"91",x"cb"),
   336 => (x"70",x"80",x"71",x"48"),
   337 => (x"02",x"bf",x"6e",x"7e"),
   338 => (x"6e",x"87",x"c8",x"c0"),
   339 => (x"66",x"c8",x"4b",x"bf"),
   340 => (x"75",x"0f",x"73",x"49"),
   341 => (x"c8",x"c0",x"02",x"9d"),
   342 => (x"dd",x"f6",x"c2",x"87"),
   343 => (x"c9",x"f3",x"49",x"bf"),
   344 => (x"e4",x"d7",x"c2",x"87"),
   345 => (x"dd",x"c0",x"02",x"bf"),
   346 => (x"c7",x"c2",x"49",x"87"),
   347 => (x"02",x"98",x"70",x"87"),
   348 => (x"c2",x"87",x"d3",x"c0"),
   349 => (x"49",x"bf",x"dd",x"f6"),
   350 => (x"c0",x"87",x"ef",x"f2"),
   351 => (x"87",x"cf",x"f4",x"49"),
   352 => (x"48",x"e4",x"d7",x"c2"),
   353 => (x"8e",x"f4",x"78",x"c0"),
   354 => (x"0e",x"87",x"e9",x"f3"),
   355 => (x"5d",x"5c",x"5b",x"5e"),
   356 => (x"4c",x"71",x"1e",x"0e"),
   357 => (x"bf",x"d9",x"f6",x"c2"),
   358 => (x"a1",x"cd",x"c1",x"49"),
   359 => (x"81",x"d1",x"c1",x"4d"),
   360 => (x"9c",x"74",x"7e",x"69"),
   361 => (x"c4",x"87",x"cf",x"02"),
   362 => (x"7b",x"74",x"4b",x"a5"),
   363 => (x"bf",x"d9",x"f6",x"c2"),
   364 => (x"87",x"c8",x"f3",x"49"),
   365 => (x"9c",x"74",x"7b",x"6e"),
   366 => (x"c0",x"87",x"c4",x"05"),
   367 => (x"c1",x"87",x"c2",x"4b"),
   368 => (x"f3",x"49",x"73",x"4b"),
   369 => (x"66",x"d4",x"87",x"c9"),
   370 => (x"49",x"87",x"c7",x"02"),
   371 => (x"4a",x"70",x"87",x"da"),
   372 => (x"4a",x"c0",x"87",x"c2"),
   373 => (x"5a",x"e8",x"d7",x"c2"),
   374 => (x"87",x"d8",x"f2",x"26"),
   375 => (x"00",x"00",x"00",x"00"),
   376 => (x"00",x"00",x"00",x"00"),
   377 => (x"00",x"00",x"00",x"00"),
   378 => (x"ff",x"4a",x"71",x"1e"),
   379 => (x"72",x"49",x"bf",x"c8"),
   380 => (x"4f",x"26",x"48",x"a1"),
   381 => (x"bf",x"c8",x"ff",x"1e"),
   382 => (x"c0",x"c0",x"c2",x"89"),
   383 => (x"a9",x"c0",x"c0",x"c0"),
   384 => (x"c0",x"87",x"c4",x"01"),
   385 => (x"c1",x"87",x"c2",x"4a"),
   386 => (x"26",x"48",x"72",x"4a"),
   387 => (x"5b",x"5e",x"0e",x"4f"),
   388 => (x"71",x"0e",x"5d",x"5c"),
   389 => (x"4c",x"d4",x"ff",x"4b"),
   390 => (x"c0",x"48",x"66",x"d0"),
   391 => (x"ff",x"49",x"d6",x"78"),
   392 => (x"c3",x"87",x"c8",x"db"),
   393 => (x"49",x"6c",x"7c",x"ff"),
   394 => (x"71",x"99",x"ff",x"c3"),
   395 => (x"f0",x"c3",x"49",x"4d"),
   396 => (x"a9",x"e0",x"c1",x"99"),
   397 => (x"c3",x"87",x"cb",x"05"),
   398 => (x"48",x"6c",x"7c",x"ff"),
   399 => (x"66",x"d0",x"98",x"c3"),
   400 => (x"ff",x"c3",x"78",x"08"),
   401 => (x"49",x"4a",x"6c",x"7c"),
   402 => (x"ff",x"c3",x"31",x"c8"),
   403 => (x"71",x"4a",x"6c",x"7c"),
   404 => (x"c8",x"49",x"72",x"b2"),
   405 => (x"7c",x"ff",x"c3",x"31"),
   406 => (x"b2",x"71",x"4a",x"6c"),
   407 => (x"31",x"c8",x"49",x"72"),
   408 => (x"6c",x"7c",x"ff",x"c3"),
   409 => (x"ff",x"b2",x"71",x"4a"),
   410 => (x"e0",x"c0",x"48",x"d0"),
   411 => (x"02",x"9b",x"73",x"78"),
   412 => (x"7b",x"72",x"87",x"c2"),
   413 => (x"4d",x"26",x"48",x"75"),
   414 => (x"4b",x"26",x"4c",x"26"),
   415 => (x"26",x"1e",x"4f",x"26"),
   416 => (x"5b",x"5e",x"0e",x"4f"),
   417 => (x"86",x"f8",x"0e",x"5c"),
   418 => (x"a6",x"c8",x"1e",x"76"),
   419 => (x"87",x"fd",x"fd",x"49"),
   420 => (x"4b",x"70",x"86",x"c4"),
   421 => (x"a8",x"c3",x"48",x"6e"),
   422 => (x"87",x"f0",x"c2",x"03"),
   423 => (x"f0",x"c3",x"4a",x"73"),
   424 => (x"aa",x"d0",x"c1",x"9a"),
   425 => (x"c1",x"87",x"c7",x"02"),
   426 => (x"c2",x"05",x"aa",x"e0"),
   427 => (x"49",x"73",x"87",x"de"),
   428 => (x"c3",x"02",x"99",x"c8"),
   429 => (x"87",x"c6",x"ff",x"87"),
   430 => (x"9c",x"c3",x"4c",x"73"),
   431 => (x"c1",x"05",x"ac",x"c2"),
   432 => (x"66",x"c4",x"87",x"c2"),
   433 => (x"71",x"31",x"c9",x"49"),
   434 => (x"4a",x"66",x"c4",x"1e"),
   435 => (x"f6",x"c2",x"92",x"d4"),
   436 => (x"81",x"72",x"49",x"e1"),
   437 => (x"87",x"fa",x"cb",x"fe"),
   438 => (x"d8",x"ff",x"49",x"d8"),
   439 => (x"c0",x"c8",x"87",x"cd"),
   440 => (x"fe",x"e4",x"c2",x"1e"),
   441 => (x"f6",x"e7",x"fd",x"49"),
   442 => (x"48",x"d0",x"ff",x"87"),
   443 => (x"c2",x"78",x"e0",x"c0"),
   444 => (x"cc",x"1e",x"fe",x"e4"),
   445 => (x"92",x"d4",x"4a",x"66"),
   446 => (x"49",x"e1",x"f6",x"c2"),
   447 => (x"ca",x"fe",x"81",x"72"),
   448 => (x"86",x"cc",x"87",x"c1"),
   449 => (x"c1",x"05",x"ac",x"c1"),
   450 => (x"66",x"c4",x"87",x"c2"),
   451 => (x"71",x"31",x"c9",x"49"),
   452 => (x"4a",x"66",x"c4",x"1e"),
   453 => (x"f6",x"c2",x"92",x"d4"),
   454 => (x"81",x"72",x"49",x"e1"),
   455 => (x"87",x"f2",x"ca",x"fe"),
   456 => (x"1e",x"fe",x"e4",x"c2"),
   457 => (x"d4",x"4a",x"66",x"c8"),
   458 => (x"e1",x"f6",x"c2",x"92"),
   459 => (x"fe",x"81",x"72",x"49"),
   460 => (x"d7",x"87",x"c1",x"c8"),
   461 => (x"f2",x"d6",x"ff",x"49"),
   462 => (x"1e",x"c0",x"c8",x"87"),
   463 => (x"49",x"fe",x"e4",x"c2"),
   464 => (x"87",x"f4",x"e5",x"fd"),
   465 => (x"d0",x"ff",x"86",x"cc"),
   466 => (x"78",x"e0",x"c0",x"48"),
   467 => (x"e7",x"fc",x"8e",x"f8"),
   468 => (x"5b",x"5e",x"0e",x"87"),
   469 => (x"1e",x"0e",x"5d",x"5c"),
   470 => (x"d4",x"ff",x"4d",x"71"),
   471 => (x"7e",x"66",x"d4",x"4c"),
   472 => (x"a8",x"b7",x"c3",x"48"),
   473 => (x"c0",x"87",x"c5",x"06"),
   474 => (x"87",x"e2",x"c1",x"48"),
   475 => (x"d8",x"fe",x"49",x"75"),
   476 => (x"1e",x"75",x"87",x"ed"),
   477 => (x"d4",x"4b",x"66",x"c4"),
   478 => (x"e1",x"f6",x"c2",x"93"),
   479 => (x"fe",x"49",x"73",x"83"),
   480 => (x"c8",x"87",x"fe",x"c1"),
   481 => (x"ff",x"4b",x"6b",x"83"),
   482 => (x"e1",x"c8",x"48",x"d0"),
   483 => (x"73",x"7c",x"dd",x"78"),
   484 => (x"99",x"ff",x"c3",x"49"),
   485 => (x"49",x"73",x"7c",x"71"),
   486 => (x"c3",x"29",x"b7",x"c8"),
   487 => (x"7c",x"71",x"99",x"ff"),
   488 => (x"b7",x"d0",x"49",x"73"),
   489 => (x"99",x"ff",x"c3",x"29"),
   490 => (x"49",x"73",x"7c",x"71"),
   491 => (x"71",x"29",x"b7",x"d8"),
   492 => (x"7c",x"7c",x"c0",x"7c"),
   493 => (x"7c",x"7c",x"7c",x"7c"),
   494 => (x"7c",x"7c",x"7c",x"7c"),
   495 => (x"e0",x"c0",x"7c",x"7c"),
   496 => (x"1e",x"66",x"c4",x"78"),
   497 => (x"d5",x"ff",x"49",x"dc"),
   498 => (x"86",x"c8",x"87",x"c6"),
   499 => (x"fa",x"26",x"48",x"73"),
   500 => (x"c2",x"1e",x"87",x"e4"),
   501 => (x"49",x"bf",x"de",x"e2"),
   502 => (x"e2",x"c2",x"b9",x"c1"),
   503 => (x"d4",x"ff",x"59",x"e2"),
   504 => (x"78",x"ff",x"c3",x"48"),
   505 => (x"c0",x"48",x"d0",x"ff"),
   506 => (x"d4",x"ff",x"78",x"e1"),
   507 => (x"c4",x"78",x"c1",x"48"),
   508 => (x"ff",x"78",x"71",x"31"),
   509 => (x"e0",x"c0",x"48",x"d0"),
   510 => (x"1e",x"4f",x"26",x"78"),
   511 => (x"a2",x"c4",x"4a",x"71"),
   512 => (x"f8",x"f5",x"c2",x"49"),
   513 => (x"69",x"78",x"6a",x"48"),
   514 => (x"c2",x"b9",x"c1",x"49"),
   515 => (x"ff",x"59",x"e2",x"e2"),
   516 => (x"d5",x"ff",x"87",x"c0"),
   517 => (x"48",x"c1",x"87",x"d4"),
   518 => (x"71",x"1e",x"4f",x"26"),
   519 => (x"49",x"a2",x"c4",x"4a"),
   520 => (x"bf",x"f8",x"f5",x"c2"),
   521 => (x"de",x"e2",x"c2",x"7a"),
   522 => (x"4f",x"26",x"79",x"bf"),
   523 => (x"9a",x"4a",x"71",x"1e"),
   524 => (x"87",x"ec",x"c0",x"02"),
   525 => (x"f4",x"f1",x"c2",x"1e"),
   526 => (x"c4",x"ff",x"fd",x"49"),
   527 => (x"70",x"86",x"c4",x"87"),
   528 => (x"87",x"dc",x"02",x"98"),
   529 => (x"1e",x"fe",x"e4",x"c2"),
   530 => (x"49",x"f4",x"f1",x"c2"),
   531 => (x"87",x"e4",x"c3",x"fe"),
   532 => (x"98",x"70",x"86",x"c4"),
   533 => (x"c2",x"87",x"c9",x"02"),
   534 => (x"fe",x"49",x"fe",x"e4"),
   535 => (x"87",x"c2",x"87",x"dd"),
   536 => (x"4f",x"26",x"48",x"c0"),
   537 => (x"9a",x"4a",x"71",x"1e"),
   538 => (x"87",x"ee",x"c0",x"02"),
   539 => (x"f4",x"f1",x"c2",x"1e"),
   540 => (x"cc",x"fe",x"fd",x"49"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"87",x"de",x"02",x"98"),
   543 => (x"49",x"fe",x"e4",x"c2"),
   544 => (x"c2",x"87",x"d7",x"fe"),
   545 => (x"c2",x"1e",x"fe",x"e4"),
   546 => (x"fe",x"49",x"f4",x"f1"),
   547 => (x"c4",x"87",x"f4",x"c3"),
   548 => (x"02",x"98",x"70",x"86"),
   549 => (x"48",x"c1",x"87",x"c4"),
   550 => (x"48",x"c0",x"87",x"c2"),
   551 => (x"00",x"00",x"4f",x"26"),
   552 => (x"73",x"1e",x"00",x"00"),
   553 => (x"c2",x"4b",x"c0",x"1e"),
   554 => (x"fd",x"49",x"d7",x"e3"),
   555 => (x"e3",x"c2",x"87",x"fe"),
   556 => (x"fe",x"49",x"bf",x"f6"),
   557 => (x"70",x"87",x"c8",x"d8"),
   558 => (x"87",x"c4",x"05",x"98"),
   559 => (x"4b",x"e3",x"e3",x"c2"),
   560 => (x"e3",x"c2",x"1e",x"c0"),
   561 => (x"fa",x"49",x"bf",x"fa"),
   562 => (x"48",x"73",x"87",x"c7"),
   563 => (x"26",x"87",x"c4",x"26"),
   564 => (x"26",x"4c",x"26",x"4d"),
   565 => (x"5a",x"4f",x"26",x"4b"),
   566 => (x"20",x"33",x"50",x"58"),
   567 => (x"43",x"20",x"20",x"20"),
   568 => (x"52",x"00",x"47",x"46"),
   569 => (x"6c",x"20",x"4d",x"4f"),
   570 => (x"69",x"64",x"61",x"6f"),
   571 => (x"66",x"20",x"67",x"6e"),
   572 => (x"65",x"6c",x"69",x"61"),
   573 => (x"28",x"fe",x"00",x"64"),
   574 => (x"29",x"0a",x"00",x"00"),
   575 => (x"58",x"5a",x"00",x"00"),
   576 => (x"20",x"20",x"33",x"50"),
   577 => (x"4f",x"52",x"20",x"20"),
   578 => (x"58",x"5a",x"00",x"4d"),
   579 => (x"20",x"20",x"33",x"50"),
   580 => (x"48",x"56",x"20",x"20"),
   581 => (x"48",x"56",x"00",x"44"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

