//-------------------------------------------------------------------------------------------------
module pll
//-------------------------------------------------------------------------------------------------
(
	input  wire clock50,
	output wire clock56,
	output wire locked
);
//-------------------------------------------------------------------------------------------------

wire ci;

IBUFG ibufg(.I(clock50), .O(ci));

PLL_BASE #
(
	.CLKIN_PERIOD  (20.000),
	.CLKFBOUT_MULT (25    ),
	.CLKOUT0_DIVIDE(11    ),
	.DIVCLK_DIVIDE ( 2    )
)
pll
(
	.RST     (1'b0  ),
	.CLKIN   (ci    ),
	.CLKFBIN (fi    ),
	.CLKFBOUT(fo    ),
	.CLKOUT0 (co    ),
	.CLKOUT1 (      ),
	.CLKOUT2 (      ),
	.CLKOUT3 (      ),
	.CLKOUT4 (      ),
	.CLKOUT5 (      ),
	.LOCKED  (locked)
);

BUFG bufg_fb(.I(fo), .O(fi));
BUFG bufg_co(.I(co), .O(clock56));

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
