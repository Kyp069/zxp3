
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e0",x"f7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e0",x"f7",x"c2"),
    14 => (x"48",x"d8",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c1",x"e6"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d4",x"02",x"99",x"71"),
    50 => (x"ff",x"48",x"12",x"87"),
    51 => (x"c4",x"78",x"08",x"d4"),
    52 => (x"c1",x"48",x"49",x"66"),
    53 => (x"58",x"a6",x"c8",x"88"),
    54 => (x"ec",x"05",x"99",x"71"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"66",x"c4",x"4a",x"71"),
    57 => (x"88",x"c1",x"48",x"49"),
    58 => (x"71",x"58",x"a6",x"c8"),
    59 => (x"87",x"d6",x"02",x"99"),
    60 => (x"c3",x"48",x"d4",x"ff"),
    61 => (x"52",x"68",x"78",x"ff"),
    62 => (x"48",x"49",x"66",x"c4"),
    63 => (x"a6",x"c8",x"88",x"c1"),
    64 => (x"05",x"99",x"71",x"58"),
    65 => (x"4f",x"26",x"87",x"ea"),
    66 => (x"ff",x"1e",x"73",x"1e"),
    67 => (x"ff",x"c3",x"4b",x"d4"),
    68 => (x"c3",x"4a",x"6b",x"7b"),
    69 => (x"49",x"6b",x"7b",x"ff"),
    70 => (x"b1",x"72",x"32",x"c8"),
    71 => (x"6b",x"7b",x"ff",x"c3"),
    72 => (x"71",x"31",x"c8",x"4a"),
    73 => (x"7b",x"ff",x"c3",x"b2"),
    74 => (x"32",x"c8",x"49",x"6b"),
    75 => (x"48",x"71",x"b1",x"72"),
    76 => (x"4d",x"26",x"87",x"c4"),
    77 => (x"4b",x"26",x"4c",x"26"),
    78 => (x"5e",x"0e",x"4f",x"26"),
    79 => (x"0e",x"5d",x"5c",x"5b"),
    80 => (x"d4",x"ff",x"4a",x"71"),
    81 => (x"c3",x"49",x"72",x"4c"),
    82 => (x"7c",x"71",x"99",x"ff"),
    83 => (x"bf",x"d8",x"e4",x"c2"),
    84 => (x"d0",x"87",x"c8",x"05"),
    85 => (x"30",x"c9",x"48",x"66"),
    86 => (x"d0",x"58",x"a6",x"d4"),
    87 => (x"29",x"d8",x"49",x"66"),
    88 => (x"71",x"99",x"ff",x"c3"),
    89 => (x"49",x"66",x"d0",x"7c"),
    90 => (x"ff",x"c3",x"29",x"d0"),
    91 => (x"d0",x"7c",x"71",x"99"),
    92 => (x"29",x"c8",x"49",x"66"),
    93 => (x"71",x"99",x"ff",x"c3"),
    94 => (x"49",x"66",x"d0",x"7c"),
    95 => (x"71",x"99",x"ff",x"c3"),
    96 => (x"d0",x"49",x"72",x"7c"),
    97 => (x"99",x"ff",x"c3",x"29"),
    98 => (x"4b",x"6c",x"7c",x"71"),
    99 => (x"4d",x"ff",x"f0",x"c9"),
   100 => (x"05",x"ab",x"ff",x"c3"),
   101 => (x"ff",x"c3",x"87",x"d0"),
   102 => (x"c1",x"4b",x"6c",x"7c"),
   103 => (x"87",x"c6",x"02",x"8d"),
   104 => (x"02",x"ab",x"ff",x"c3"),
   105 => (x"48",x"73",x"87",x"f0"),
   106 => (x"1e",x"87",x"c7",x"fe"),
   107 => (x"d4",x"ff",x"49",x"c0"),
   108 => (x"78",x"ff",x"c3",x"48"),
   109 => (x"c8",x"c3",x"81",x"c1"),
   110 => (x"f1",x"04",x"a9",x"b7"),
   111 => (x"1e",x"4f",x"26",x"87"),
   112 => (x"87",x"e7",x"1e",x"73"),
   113 => (x"4b",x"df",x"f8",x"c4"),
   114 => (x"ff",x"c0",x"1e",x"c0"),
   115 => (x"49",x"f7",x"c1",x"f0"),
   116 => (x"c4",x"87",x"e7",x"fd"),
   117 => (x"05",x"a8",x"c1",x"86"),
   118 => (x"ff",x"87",x"ea",x"c0"),
   119 => (x"ff",x"c3",x"48",x"d4"),
   120 => (x"c0",x"c0",x"c1",x"78"),
   121 => (x"1e",x"c0",x"c0",x"c0"),
   122 => (x"c1",x"f0",x"e1",x"c0"),
   123 => (x"c9",x"fd",x"49",x"e9"),
   124 => (x"70",x"86",x"c4",x"87"),
   125 => (x"87",x"ca",x"05",x"98"),
   126 => (x"c3",x"48",x"d4",x"ff"),
   127 => (x"48",x"c1",x"78",x"ff"),
   128 => (x"e6",x"fe",x"87",x"cb"),
   129 => (x"05",x"8b",x"c1",x"87"),
   130 => (x"c0",x"87",x"fd",x"fe"),
   131 => (x"87",x"e6",x"fc",x"48"),
   132 => (x"ff",x"1e",x"73",x"1e"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"c0",x"4b",x"d3",x"78"),
   135 => (x"f0",x"ff",x"c0",x"1e"),
   136 => (x"fc",x"49",x"c1",x"c1"),
   137 => (x"86",x"c4",x"87",x"d4"),
   138 => (x"ca",x"05",x"98",x"70"),
   139 => (x"48",x"d4",x"ff",x"87"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"fd",x"87",x"cb",x"48"),
   142 => (x"8b",x"c1",x"87",x"f1"),
   143 => (x"87",x"db",x"ff",x"05"),
   144 => (x"f1",x"fb",x"48",x"c0"),
   145 => (x"5b",x"5e",x"0e",x"87"),
   146 => (x"d4",x"ff",x"0e",x"5c"),
   147 => (x"87",x"db",x"fd",x"4c"),
   148 => (x"c0",x"1e",x"ea",x"c6"),
   149 => (x"c8",x"c1",x"f0",x"e1"),
   150 => (x"87",x"de",x"fb",x"49"),
   151 => (x"a8",x"c1",x"86",x"c4"),
   152 => (x"fe",x"87",x"c8",x"02"),
   153 => (x"48",x"c0",x"87",x"ea"),
   154 => (x"fa",x"87",x"e2",x"c1"),
   155 => (x"49",x"70",x"87",x"da"),
   156 => (x"99",x"ff",x"ff",x"cf"),
   157 => (x"02",x"a9",x"ea",x"c6"),
   158 => (x"d3",x"fe",x"87",x"c8"),
   159 => (x"c1",x"48",x"c0",x"87"),
   160 => (x"ff",x"c3",x"87",x"cb"),
   161 => (x"4b",x"f1",x"c0",x"7c"),
   162 => (x"70",x"87",x"f4",x"fc"),
   163 => (x"eb",x"c0",x"02",x"98"),
   164 => (x"c0",x"1e",x"c0",x"87"),
   165 => (x"fa",x"c1",x"f0",x"ff"),
   166 => (x"87",x"de",x"fa",x"49"),
   167 => (x"98",x"70",x"86",x"c4"),
   168 => (x"c3",x"87",x"d9",x"05"),
   169 => (x"49",x"6c",x"7c",x"ff"),
   170 => (x"7c",x"7c",x"ff",x"c3"),
   171 => (x"c0",x"c1",x"7c",x"7c"),
   172 => (x"87",x"c4",x"02",x"99"),
   173 => (x"87",x"d5",x"48",x"c1"),
   174 => (x"87",x"d1",x"48",x"c0"),
   175 => (x"c4",x"05",x"ab",x"c2"),
   176 => (x"c8",x"48",x"c0",x"87"),
   177 => (x"05",x"8b",x"c1",x"87"),
   178 => (x"c0",x"87",x"fd",x"fe"),
   179 => (x"87",x"e4",x"f9",x"48"),
   180 => (x"c2",x"1e",x"73",x"1e"),
   181 => (x"c1",x"48",x"d8",x"e4"),
   182 => (x"ff",x"4b",x"c7",x"78"),
   183 => (x"78",x"c2",x"48",x"d0"),
   184 => (x"ff",x"87",x"c8",x"fb"),
   185 => (x"78",x"c3",x"48",x"d0"),
   186 => (x"e5",x"c0",x"1e",x"c0"),
   187 => (x"49",x"c0",x"c1",x"d0"),
   188 => (x"c4",x"87",x"c7",x"f9"),
   189 => (x"05",x"a8",x"c1",x"86"),
   190 => (x"c2",x"4b",x"87",x"c1"),
   191 => (x"87",x"c5",x"05",x"ab"),
   192 => (x"f9",x"c0",x"48",x"c0"),
   193 => (x"05",x"8b",x"c1",x"87"),
   194 => (x"fc",x"87",x"d0",x"ff"),
   195 => (x"e4",x"c2",x"87",x"f7"),
   196 => (x"98",x"70",x"58",x"dc"),
   197 => (x"c1",x"87",x"cd",x"05"),
   198 => (x"f0",x"ff",x"c0",x"1e"),
   199 => (x"f8",x"49",x"d0",x"c1"),
   200 => (x"86",x"c4",x"87",x"d8"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"de",x"c4",x"78",x"ff"),
   203 => (x"e0",x"e4",x"c2",x"87"),
   204 => (x"48",x"d0",x"ff",x"58"),
   205 => (x"d4",x"ff",x"78",x"c2"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"f5",x"f7",x"48",x"c1"),
   208 => (x"5b",x"5e",x"0e",x"87"),
   209 => (x"71",x"0e",x"5d",x"5c"),
   210 => (x"4d",x"ff",x"c3",x"4a"),
   211 => (x"75",x"4c",x"d4",x"ff"),
   212 => (x"48",x"d0",x"ff",x"7c"),
   213 => (x"75",x"78",x"c3",x"c4"),
   214 => (x"c0",x"1e",x"72",x"7c"),
   215 => (x"d8",x"c1",x"f0",x"ff"),
   216 => (x"87",x"d6",x"f7",x"49"),
   217 => (x"98",x"70",x"86",x"c4"),
   218 => (x"c1",x"87",x"c5",x"02"),
   219 => (x"87",x"f0",x"c0",x"48"),
   220 => (x"fe",x"c3",x"7c",x"75"),
   221 => (x"1e",x"c0",x"c8",x"7c"),
   222 => (x"f4",x"49",x"66",x"d4"),
   223 => (x"86",x"c4",x"87",x"fa"),
   224 => (x"7c",x"75",x"7c",x"75"),
   225 => (x"da",x"d8",x"7c",x"75"),
   226 => (x"7c",x"75",x"4b",x"e0"),
   227 => (x"05",x"99",x"49",x"6c"),
   228 => (x"8b",x"c1",x"87",x"c5"),
   229 => (x"75",x"87",x"f3",x"05"),
   230 => (x"48",x"d0",x"ff",x"7c"),
   231 => (x"48",x"c0",x"78",x"c2"),
   232 => (x"0e",x"87",x"cf",x"f6"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"4b",x"71",x"0e"),
   235 => (x"cd",x"ee",x"c5",x"4c"),
   236 => (x"d4",x"ff",x"4a",x"df"),
   237 => (x"78",x"ff",x"c3",x"48"),
   238 => (x"fe",x"c3",x"49",x"68"),
   239 => (x"fd",x"c0",x"05",x"a9"),
   240 => (x"73",x"4d",x"70",x"87"),
   241 => (x"87",x"cc",x"02",x"9b"),
   242 => (x"73",x"1e",x"66",x"d0"),
   243 => (x"87",x"cf",x"f4",x"49"),
   244 => (x"87",x"d6",x"86",x"c4"),
   245 => (x"c4",x"48",x"d0",x"ff"),
   246 => (x"ff",x"c3",x"78",x"d1"),
   247 => (x"48",x"66",x"d0",x"7d"),
   248 => (x"a6",x"d4",x"88",x"c1"),
   249 => (x"05",x"98",x"70",x"58"),
   250 => (x"d4",x"ff",x"87",x"f0"),
   251 => (x"78",x"ff",x"c3",x"48"),
   252 => (x"05",x"9b",x"73",x"78"),
   253 => (x"d0",x"ff",x"87",x"c5"),
   254 => (x"c1",x"78",x"d0",x"48"),
   255 => (x"8a",x"c1",x"4c",x"4a"),
   256 => (x"87",x"ee",x"fe",x"05"),
   257 => (x"e9",x"f4",x"48",x"74"),
   258 => (x"1e",x"73",x"1e",x"87"),
   259 => (x"4b",x"c0",x"4a",x"71"),
   260 => (x"c3",x"48",x"d4",x"ff"),
   261 => (x"d0",x"ff",x"78",x"ff"),
   262 => (x"78",x"c3",x"c4",x"48"),
   263 => (x"c3",x"48",x"d4",x"ff"),
   264 => (x"1e",x"72",x"78",x"ff"),
   265 => (x"c1",x"f0",x"ff",x"c0"),
   266 => (x"cd",x"f4",x"49",x"d1"),
   267 => (x"70",x"86",x"c4",x"87"),
   268 => (x"87",x"d2",x"05",x"98"),
   269 => (x"cc",x"1e",x"c0",x"c8"),
   270 => (x"e6",x"fd",x"49",x"66"),
   271 => (x"70",x"86",x"c4",x"87"),
   272 => (x"48",x"d0",x"ff",x"4b"),
   273 => (x"48",x"73",x"78",x"c2"),
   274 => (x"0e",x"87",x"eb",x"f3"),
   275 => (x"5d",x"5c",x"5b",x"5e"),
   276 => (x"c0",x"1e",x"c0",x"0e"),
   277 => (x"c9",x"c1",x"f0",x"ff"),
   278 => (x"87",x"de",x"f3",x"49"),
   279 => (x"e4",x"c2",x"1e",x"d2"),
   280 => (x"fe",x"fc",x"49",x"e0"),
   281 => (x"c0",x"86",x"c8",x"87"),
   282 => (x"d2",x"84",x"c1",x"4c"),
   283 => (x"f8",x"04",x"ac",x"b7"),
   284 => (x"e0",x"e4",x"c2",x"87"),
   285 => (x"c3",x"49",x"bf",x"97"),
   286 => (x"c0",x"c1",x"99",x"c0"),
   287 => (x"e7",x"c0",x"05",x"a9"),
   288 => (x"e7",x"e4",x"c2",x"87"),
   289 => (x"d0",x"49",x"bf",x"97"),
   290 => (x"e8",x"e4",x"c2",x"31"),
   291 => (x"c8",x"4a",x"bf",x"97"),
   292 => (x"c2",x"b1",x"72",x"32"),
   293 => (x"bf",x"97",x"e9",x"e4"),
   294 => (x"4c",x"71",x"b1",x"4a"),
   295 => (x"ff",x"ff",x"ff",x"cf"),
   296 => (x"ca",x"84",x"c1",x"9c"),
   297 => (x"87",x"e7",x"c1",x"34"),
   298 => (x"97",x"e9",x"e4",x"c2"),
   299 => (x"31",x"c1",x"49",x"bf"),
   300 => (x"e4",x"c2",x"99",x"c6"),
   301 => (x"4a",x"bf",x"97",x"ea"),
   302 => (x"72",x"2a",x"b7",x"c7"),
   303 => (x"e5",x"e4",x"c2",x"b1"),
   304 => (x"4d",x"4a",x"bf",x"97"),
   305 => (x"e4",x"c2",x"9d",x"cf"),
   306 => (x"4a",x"bf",x"97",x"e6"),
   307 => (x"32",x"ca",x"9a",x"c3"),
   308 => (x"97",x"e7",x"e4",x"c2"),
   309 => (x"33",x"c2",x"4b",x"bf"),
   310 => (x"e4",x"c2",x"b2",x"73"),
   311 => (x"4b",x"bf",x"97",x"e8"),
   312 => (x"c6",x"9b",x"c0",x"c3"),
   313 => (x"b2",x"73",x"2b",x"b7"),
   314 => (x"48",x"c1",x"81",x"c2"),
   315 => (x"49",x"70",x"30",x"71"),
   316 => (x"30",x"75",x"48",x"c1"),
   317 => (x"4c",x"72",x"4d",x"70"),
   318 => (x"94",x"71",x"84",x"c1"),
   319 => (x"ad",x"b7",x"c0",x"c8"),
   320 => (x"c1",x"87",x"cc",x"06"),
   321 => (x"c8",x"2d",x"b7",x"34"),
   322 => (x"01",x"ad",x"b7",x"c0"),
   323 => (x"74",x"87",x"f4",x"ff"),
   324 => (x"87",x"de",x"f0",x"48"),
   325 => (x"5c",x"5b",x"5e",x"0e"),
   326 => (x"86",x"f8",x"0e",x"5d"),
   327 => (x"48",x"c6",x"ed",x"c2"),
   328 => (x"e4",x"c2",x"78",x"c0"),
   329 => (x"49",x"c0",x"1e",x"fe"),
   330 => (x"c4",x"87",x"de",x"fb"),
   331 => (x"05",x"98",x"70",x"86"),
   332 => (x"48",x"c0",x"87",x"c5"),
   333 => (x"c0",x"87",x"ce",x"c9"),
   334 => (x"c0",x"7e",x"c1",x"4d"),
   335 => (x"49",x"bf",x"ed",x"f2"),
   336 => (x"4a",x"f4",x"e5",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"e0"),
   339 => (x"c0",x"87",x"c2",x"05"),
   340 => (x"e9",x"f2",x"c0",x"7e"),
   341 => (x"e6",x"c2",x"49",x"bf"),
   342 => (x"c8",x"71",x"4a",x"d0"),
   343 => (x"87",x"ca",x"ec",x"4b"),
   344 => (x"c2",x"05",x"98",x"70"),
   345 => (x"6e",x"7e",x"c0",x"87"),
   346 => (x"87",x"fd",x"c0",x"02"),
   347 => (x"bf",x"c4",x"ec",x"c2"),
   348 => (x"fc",x"ec",x"c2",x"4d"),
   349 => (x"48",x"7e",x"bf",x"9f"),
   350 => (x"a8",x"ea",x"d6",x"c5"),
   351 => (x"c2",x"87",x"c7",x"05"),
   352 => (x"4d",x"bf",x"c4",x"ec"),
   353 => (x"48",x"6e",x"87",x"ce"),
   354 => (x"a8",x"d5",x"e9",x"ca"),
   355 => (x"c0",x"87",x"c5",x"02"),
   356 => (x"87",x"f1",x"c7",x"48"),
   357 => (x"1e",x"fe",x"e4",x"c2"),
   358 => (x"ec",x"f9",x"49",x"75"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"dc",x"c7",x"48",x"c0"),
   362 => (x"e9",x"f2",x"c0",x"87"),
   363 => (x"e6",x"c2",x"49",x"bf"),
   364 => (x"c8",x"71",x"4a",x"d0"),
   365 => (x"87",x"f2",x"ea",x"4b"),
   366 => (x"c8",x"05",x"98",x"70"),
   367 => (x"c6",x"ed",x"c2",x"87"),
   368 => (x"da",x"78",x"c1",x"48"),
   369 => (x"ed",x"f2",x"c0",x"87"),
   370 => (x"e5",x"c2",x"49",x"bf"),
   371 => (x"c8",x"71",x"4a",x"f4"),
   372 => (x"87",x"d6",x"ea",x"4b"),
   373 => (x"c0",x"02",x"98",x"70"),
   374 => (x"48",x"c0",x"87",x"c5"),
   375 => (x"c2",x"87",x"e6",x"c6"),
   376 => (x"bf",x"97",x"fc",x"ec"),
   377 => (x"a9",x"d5",x"c1",x"49"),
   378 => (x"87",x"cd",x"c0",x"05"),
   379 => (x"97",x"fd",x"ec",x"c2"),
   380 => (x"ea",x"c2",x"49",x"bf"),
   381 => (x"c5",x"c0",x"02",x"a9"),
   382 => (x"c6",x"48",x"c0",x"87"),
   383 => (x"e4",x"c2",x"87",x"c7"),
   384 => (x"7e",x"bf",x"97",x"fe"),
   385 => (x"a8",x"e9",x"c3",x"48"),
   386 => (x"87",x"ce",x"c0",x"02"),
   387 => (x"eb",x"c3",x"48",x"6e"),
   388 => (x"c5",x"c0",x"02",x"a8"),
   389 => (x"c5",x"48",x"c0",x"87"),
   390 => (x"e5",x"c2",x"87",x"eb"),
   391 => (x"49",x"bf",x"97",x"c9"),
   392 => (x"cc",x"c0",x"05",x"99"),
   393 => (x"ca",x"e5",x"c2",x"87"),
   394 => (x"c2",x"49",x"bf",x"97"),
   395 => (x"c5",x"c0",x"02",x"a9"),
   396 => (x"c5",x"48",x"c0",x"87"),
   397 => (x"e5",x"c2",x"87",x"cf"),
   398 => (x"48",x"bf",x"97",x"cb"),
   399 => (x"58",x"c2",x"ed",x"c2"),
   400 => (x"c1",x"48",x"4c",x"70"),
   401 => (x"c6",x"ed",x"c2",x"88"),
   402 => (x"cc",x"e5",x"c2",x"58"),
   403 => (x"75",x"49",x"bf",x"97"),
   404 => (x"cd",x"e5",x"c2",x"81"),
   405 => (x"c8",x"4a",x"bf",x"97"),
   406 => (x"7e",x"a1",x"72",x"32"),
   407 => (x"48",x"d3",x"f1",x"c2"),
   408 => (x"e5",x"c2",x"78",x"6e"),
   409 => (x"48",x"bf",x"97",x"ce"),
   410 => (x"c2",x"58",x"a6",x"c8"),
   411 => (x"02",x"bf",x"c6",x"ed"),
   412 => (x"c0",x"87",x"d4",x"c2"),
   413 => (x"49",x"bf",x"e9",x"f2"),
   414 => (x"4a",x"d0",x"e6",x"c2"),
   415 => (x"e7",x"4b",x"c8",x"71"),
   416 => (x"98",x"70",x"87",x"e8"),
   417 => (x"87",x"c5",x"c0",x"02"),
   418 => (x"f8",x"c3",x"48",x"c0"),
   419 => (x"fe",x"ec",x"c2",x"87"),
   420 => (x"f1",x"c2",x"4c",x"bf"),
   421 => (x"e5",x"c2",x"5c",x"e7"),
   422 => (x"49",x"bf",x"97",x"e3"),
   423 => (x"e5",x"c2",x"31",x"c8"),
   424 => (x"4a",x"bf",x"97",x"e2"),
   425 => (x"e5",x"c2",x"49",x"a1"),
   426 => (x"4a",x"bf",x"97",x"e4"),
   427 => (x"a1",x"72",x"32",x"d0"),
   428 => (x"e5",x"e5",x"c2",x"49"),
   429 => (x"d8",x"4a",x"bf",x"97"),
   430 => (x"49",x"a1",x"72",x"32"),
   431 => (x"c2",x"91",x"66",x"c4"),
   432 => (x"81",x"bf",x"d3",x"f1"),
   433 => (x"59",x"db",x"f1",x"c2"),
   434 => (x"97",x"eb",x"e5",x"c2"),
   435 => (x"32",x"c8",x"4a",x"bf"),
   436 => (x"97",x"ea",x"e5",x"c2"),
   437 => (x"4a",x"a2",x"4b",x"bf"),
   438 => (x"97",x"ec",x"e5",x"c2"),
   439 => (x"33",x"d0",x"4b",x"bf"),
   440 => (x"c2",x"4a",x"a2",x"73"),
   441 => (x"bf",x"97",x"ed",x"e5"),
   442 => (x"d8",x"9b",x"cf",x"4b"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"5a",x"df",x"f1",x"c2"),
   445 => (x"bf",x"db",x"f1",x"c2"),
   446 => (x"74",x"8a",x"c2",x"4a"),
   447 => (x"df",x"f1",x"c2",x"92"),
   448 => (x"78",x"a1",x"72",x"48"),
   449 => (x"c2",x"87",x"ca",x"c1"),
   450 => (x"bf",x"97",x"d0",x"e5"),
   451 => (x"c2",x"31",x"c8",x"49"),
   452 => (x"bf",x"97",x"cf",x"e5"),
   453 => (x"c2",x"49",x"a1",x"4a"),
   454 => (x"c2",x"59",x"ce",x"ed"),
   455 => (x"49",x"bf",x"ca",x"ed"),
   456 => (x"ff",x"c7",x"31",x"c5"),
   457 => (x"c2",x"29",x"c9",x"81"),
   458 => (x"c2",x"59",x"e7",x"f1"),
   459 => (x"bf",x"97",x"d5",x"e5"),
   460 => (x"c2",x"32",x"c8",x"4a"),
   461 => (x"bf",x"97",x"d4",x"e5"),
   462 => (x"c4",x"4a",x"a2",x"4b"),
   463 => (x"82",x"6e",x"92",x"66"),
   464 => (x"5a",x"e3",x"f1",x"c2"),
   465 => (x"48",x"db",x"f1",x"c2"),
   466 => (x"f1",x"c2",x"78",x"c0"),
   467 => (x"a1",x"72",x"48",x"d7"),
   468 => (x"e7",x"f1",x"c2",x"78"),
   469 => (x"db",x"f1",x"c2",x"48"),
   470 => (x"f1",x"c2",x"78",x"bf"),
   471 => (x"f1",x"c2",x"48",x"eb"),
   472 => (x"c2",x"78",x"bf",x"df"),
   473 => (x"02",x"bf",x"c6",x"ed"),
   474 => (x"74",x"87",x"c9",x"c0"),
   475 => (x"70",x"30",x"c4",x"48"),
   476 => (x"87",x"c9",x"c0",x"7e"),
   477 => (x"bf",x"e3",x"f1",x"c2"),
   478 => (x"70",x"30",x"c4",x"48"),
   479 => (x"ca",x"ed",x"c2",x"7e"),
   480 => (x"c1",x"78",x"6e",x"48"),
   481 => (x"26",x"8e",x"f8",x"48"),
   482 => (x"26",x"4c",x"26",x"4d"),
   483 => (x"0e",x"4f",x"26",x"4b"),
   484 => (x"5d",x"5c",x"5b",x"5e"),
   485 => (x"c2",x"4a",x"71",x"0e"),
   486 => (x"02",x"bf",x"c6",x"ed"),
   487 => (x"4b",x"72",x"87",x"cb"),
   488 => (x"4c",x"72",x"2b",x"c7"),
   489 => (x"c9",x"9c",x"ff",x"c1"),
   490 => (x"c8",x"4b",x"72",x"87"),
   491 => (x"c3",x"4c",x"72",x"2b"),
   492 => (x"f1",x"c2",x"9c",x"ff"),
   493 => (x"c0",x"83",x"bf",x"d3"),
   494 => (x"ab",x"bf",x"e5",x"f2"),
   495 => (x"c0",x"87",x"d9",x"02"),
   496 => (x"c2",x"5b",x"e9",x"f2"),
   497 => (x"73",x"1e",x"fe",x"e4"),
   498 => (x"87",x"fd",x"f0",x"49"),
   499 => (x"98",x"70",x"86",x"c4"),
   500 => (x"c0",x"87",x"c5",x"05"),
   501 => (x"87",x"e6",x"c0",x"48"),
   502 => (x"bf",x"c6",x"ed",x"c2"),
   503 => (x"74",x"87",x"d2",x"02"),
   504 => (x"c2",x"91",x"c4",x"49"),
   505 => (x"69",x"81",x"fe",x"e4"),
   506 => (x"ff",x"ff",x"cf",x"4d"),
   507 => (x"cb",x"9d",x"ff",x"ff"),
   508 => (x"c2",x"49",x"74",x"87"),
   509 => (x"fe",x"e4",x"c2",x"91"),
   510 => (x"4d",x"69",x"9f",x"81"),
   511 => (x"c6",x"fe",x"48",x"75"),
   512 => (x"5b",x"5e",x"0e",x"87"),
   513 => (x"f8",x"0e",x"5d",x"5c"),
   514 => (x"9c",x"4c",x"71",x"86"),
   515 => (x"c0",x"87",x"c5",x"05"),
   516 => (x"87",x"c1",x"c3",x"48"),
   517 => (x"6e",x"7e",x"a4",x"c8"),
   518 => (x"d8",x"78",x"c0",x"48"),
   519 => (x"87",x"c7",x"02",x"66"),
   520 => (x"bf",x"97",x"66",x"d8"),
   521 => (x"c0",x"87",x"c5",x"05"),
   522 => (x"87",x"e9",x"c2",x"48"),
   523 => (x"49",x"c1",x"1e",x"c0"),
   524 => (x"c4",x"87",x"d7",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"ce",x"ed",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c9"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ee"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"d5",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"c6",x"ed"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ed"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"c2",x"ed",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fc",x"f9"),
   581 => (x"fe",x"ec",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"c2",x"ed",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d3",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"d7",x"f1",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"fe",x"ec",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"c2",x"ed",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"e9",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d6",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c8",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"d7",x"f1",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"fe",x"ec",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"c2",x"ed",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"e9"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"ff"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f9"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"d4",x"4b",x"71",x"1e"),
   631 => (x"9b",x"73",x"4d",x"66"),
   632 => (x"87",x"cc",x"c1",x"02"),
   633 => (x"69",x"49",x"a3",x"c8"),
   634 => (x"87",x"c4",x"c1",x"02"),
   635 => (x"c2",x"4c",x"a3",x"d0"),
   636 => (x"49",x"bf",x"c2",x"ed"),
   637 => (x"4a",x"6c",x"b9",x"ff"),
   638 => (x"66",x"d4",x"7e",x"99"),
   639 => (x"87",x"cd",x"06",x"a9"),
   640 => (x"cc",x"7c",x"7b",x"c0"),
   641 => (x"a3",x"c4",x"4a",x"a3"),
   642 => (x"ca",x"79",x"6a",x"49"),
   643 => (x"f8",x"49",x"72",x"87"),
   644 => (x"66",x"d4",x"99",x"c0"),
   645 => (x"75",x"8d",x"71",x"4d"),
   646 => (x"71",x"29",x"c9",x"49"),
   647 => (x"fa",x"49",x"73",x"1e"),
   648 => (x"e4",x"c2",x"87",x"f8"),
   649 => (x"49",x"73",x"1e",x"fe"),
   650 => (x"c8",x"87",x"c9",x"fc"),
   651 => (x"7c",x"66",x"d4",x"86"),
   652 => (x"87",x"d3",x"f5",x"26"),
   653 => (x"71",x"1e",x"73",x"1e"),
   654 => (x"c0",x"02",x"9b",x"4b"),
   655 => (x"f1",x"c2",x"87",x"e4"),
   656 => (x"4a",x"73",x"5b",x"eb"),
   657 => (x"ec",x"c2",x"8a",x"c2"),
   658 => (x"92",x"49",x"bf",x"fe"),
   659 => (x"bf",x"d7",x"f1",x"c2"),
   660 => (x"c2",x"80",x"72",x"48"),
   661 => (x"71",x"58",x"ef",x"f1"),
   662 => (x"c2",x"30",x"c4",x"48"),
   663 => (x"c0",x"58",x"ce",x"ed"),
   664 => (x"f1",x"c2",x"87",x"ed"),
   665 => (x"f1",x"c2",x"48",x"e7"),
   666 => (x"c2",x"78",x"bf",x"db"),
   667 => (x"c2",x"48",x"eb",x"f1"),
   668 => (x"78",x"bf",x"df",x"f1"),
   669 => (x"bf",x"c6",x"ed",x"c2"),
   670 => (x"c2",x"87",x"c9",x"02"),
   671 => (x"49",x"bf",x"fe",x"ec"),
   672 => (x"87",x"c7",x"31",x"c4"),
   673 => (x"bf",x"e3",x"f1",x"c2"),
   674 => (x"c2",x"31",x"c4",x"49"),
   675 => (x"f3",x"59",x"ce",x"ed"),
   676 => (x"5e",x"0e",x"87",x"f9"),
   677 => (x"71",x"0e",x"5c",x"5b"),
   678 => (x"72",x"4b",x"c0",x"4a"),
   679 => (x"e1",x"c0",x"02",x"9a"),
   680 => (x"49",x"a2",x"da",x"87"),
   681 => (x"c2",x"4b",x"69",x"9f"),
   682 => (x"02",x"bf",x"c6",x"ed"),
   683 => (x"a2",x"d4",x"87",x"cf"),
   684 => (x"49",x"69",x"9f",x"49"),
   685 => (x"ff",x"ff",x"c0",x"4c"),
   686 => (x"c2",x"34",x"d0",x"9c"),
   687 => (x"74",x"4c",x"c0",x"87"),
   688 => (x"49",x"73",x"b3",x"49"),
   689 => (x"f2",x"87",x"ed",x"fd"),
   690 => (x"5e",x"0e",x"87",x"ff"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4a",x"71",x"86",x"f4"),
   693 => (x"9a",x"72",x"7e",x"c0"),
   694 => (x"c2",x"87",x"d8",x"02"),
   695 => (x"c0",x"48",x"fa",x"e4"),
   696 => (x"f2",x"e4",x"c2",x"78"),
   697 => (x"eb",x"f1",x"c2",x"48"),
   698 => (x"e4",x"c2",x"78",x"bf"),
   699 => (x"f1",x"c2",x"48",x"f6"),
   700 => (x"c2",x"78",x"bf",x"e7"),
   701 => (x"c0",x"48",x"db",x"ed"),
   702 => (x"ca",x"ed",x"c2",x"50"),
   703 => (x"e4",x"c2",x"49",x"bf"),
   704 => (x"71",x"4a",x"bf",x"fa"),
   705 => (x"c9",x"c4",x"03",x"aa"),
   706 => (x"cf",x"49",x"72",x"87"),
   707 => (x"e9",x"c0",x"05",x"99"),
   708 => (x"e5",x"f2",x"c0",x"87"),
   709 => (x"f2",x"e4",x"c2",x"48"),
   710 => (x"e4",x"c2",x"78",x"bf"),
   711 => (x"e4",x"c2",x"1e",x"fe"),
   712 => (x"c2",x"49",x"bf",x"f2"),
   713 => (x"c1",x"48",x"f2",x"e4"),
   714 => (x"e3",x"71",x"78",x"a1"),
   715 => (x"86",x"c4",x"87",x"db"),
   716 => (x"48",x"e1",x"f2",x"c0"),
   717 => (x"78",x"fe",x"e4",x"c2"),
   718 => (x"f2",x"c0",x"87",x"cc"),
   719 => (x"c0",x"48",x"bf",x"e1"),
   720 => (x"f2",x"c0",x"80",x"e0"),
   721 => (x"e4",x"c2",x"58",x"e5"),
   722 => (x"c1",x"48",x"bf",x"fa"),
   723 => (x"fe",x"e4",x"c2",x"80"),
   724 => (x"0c",x"a1",x"27",x"58"),
   725 => (x"97",x"bf",x"00",x"00"),
   726 => (x"02",x"9d",x"4d",x"bf"),
   727 => (x"c3",x"87",x"e3",x"c2"),
   728 => (x"c2",x"02",x"ad",x"e5"),
   729 => (x"f2",x"c0",x"87",x"dc"),
   730 => (x"cb",x"4b",x"bf",x"e1"),
   731 => (x"4c",x"11",x"49",x"a3"),
   732 => (x"c1",x"05",x"ac",x"cf"),
   733 => (x"49",x"75",x"87",x"d2"),
   734 => (x"89",x"c1",x"99",x"df"),
   735 => (x"ed",x"c2",x"91",x"cd"),
   736 => (x"a3",x"c1",x"81",x"ce"),
   737 => (x"c3",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"c5"),
   740 => (x"4a",x"a3",x"c7",x"51"),
   741 => (x"a3",x"c9",x"51",x"12"),
   742 => (x"ce",x"51",x"12",x"4a"),
   743 => (x"51",x"12",x"4a",x"a3"),
   744 => (x"12",x"4a",x"a3",x"d0"),
   745 => (x"4a",x"a3",x"d2",x"51"),
   746 => (x"a3",x"d4",x"51",x"12"),
   747 => (x"d6",x"51",x"12",x"4a"),
   748 => (x"51",x"12",x"4a",x"a3"),
   749 => (x"12",x"4a",x"a3",x"d8"),
   750 => (x"4a",x"a3",x"dc",x"51"),
   751 => (x"a3",x"de",x"51",x"12"),
   752 => (x"c1",x"51",x"12",x"4a"),
   753 => (x"87",x"fa",x"c0",x"7e"),
   754 => (x"99",x"c8",x"49",x"74"),
   755 => (x"87",x"eb",x"c0",x"05"),
   756 => (x"99",x"d0",x"49",x"74"),
   757 => (x"dc",x"87",x"d1",x"05"),
   758 => (x"cb",x"c0",x"02",x"66"),
   759 => (x"dc",x"49",x"73",x"87"),
   760 => (x"98",x"70",x"0f",x"66"),
   761 => (x"87",x"d3",x"c0",x"02"),
   762 => (x"c6",x"c0",x"05",x"6e"),
   763 => (x"ce",x"ed",x"c2",x"87"),
   764 => (x"c0",x"50",x"c0",x"48"),
   765 => (x"48",x"bf",x"e1",x"f2"),
   766 => (x"c2",x"87",x"e1",x"c2"),
   767 => (x"c0",x"48",x"db",x"ed"),
   768 => (x"ed",x"c2",x"7e",x"50"),
   769 => (x"c2",x"49",x"bf",x"ca"),
   770 => (x"4a",x"bf",x"fa",x"e4"),
   771 => (x"fb",x"04",x"aa",x"71"),
   772 => (x"f1",x"c2",x"87",x"f7"),
   773 => (x"c0",x"05",x"bf",x"eb"),
   774 => (x"ed",x"c2",x"87",x"c8"),
   775 => (x"c1",x"02",x"bf",x"c6"),
   776 => (x"e4",x"c2",x"87",x"f8"),
   777 => (x"ed",x"49",x"bf",x"f6"),
   778 => (x"49",x"70",x"87",x"e5"),
   779 => (x"59",x"fa",x"e4",x"c2"),
   780 => (x"c2",x"48",x"a6",x"c4"),
   781 => (x"78",x"bf",x"f6",x"e4"),
   782 => (x"bf",x"c6",x"ed",x"c2"),
   783 => (x"87",x"d8",x"c0",x"02"),
   784 => (x"cf",x"49",x"66",x"c4"),
   785 => (x"f8",x"ff",x"ff",x"ff"),
   786 => (x"c0",x"02",x"a9",x"99"),
   787 => (x"4c",x"c0",x"87",x"c5"),
   788 => (x"c1",x"87",x"e1",x"c0"),
   789 => (x"87",x"dc",x"c0",x"4c"),
   790 => (x"cf",x"49",x"66",x"c4"),
   791 => (x"a9",x"99",x"f8",x"ff"),
   792 => (x"87",x"c8",x"c0",x"02"),
   793 => (x"c0",x"48",x"a6",x"c8"),
   794 => (x"87",x"c5",x"c0",x"78"),
   795 => (x"c1",x"48",x"a6",x"c8"),
   796 => (x"4c",x"66",x"c8",x"78"),
   797 => (x"c0",x"05",x"9c",x"74"),
   798 => (x"66",x"c4",x"87",x"e0"),
   799 => (x"c2",x"89",x"c2",x"49"),
   800 => (x"4a",x"bf",x"fe",x"ec"),
   801 => (x"d7",x"f1",x"c2",x"91"),
   802 => (x"e4",x"c2",x"4a",x"bf"),
   803 => (x"a1",x"72",x"48",x"f2"),
   804 => (x"fa",x"e4",x"c2",x"78"),
   805 => (x"f9",x"78",x"c0",x"48"),
   806 => (x"48",x"c0",x"87",x"df"),
   807 => (x"e6",x"eb",x"8e",x"f4"),
   808 => (x"00",x"00",x"00",x"87"),
   809 => (x"ff",x"ff",x"ff",x"00"),
   810 => (x"00",x"0c",x"b1",x"ff"),
   811 => (x"00",x"0c",x"ba",x"00"),
   812 => (x"54",x"41",x"46",x"00"),
   813 => (x"20",x"20",x"32",x"33"),
   814 => (x"41",x"46",x"00",x"20"),
   815 => (x"20",x"36",x"31",x"54"),
   816 => (x"1e",x"00",x"20",x"20"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"48",x"68",x"78",x"ff"),
   819 => (x"ff",x"1e",x"4f",x"26"),
   820 => (x"ff",x"c3",x"48",x"d4"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"ff",x"78",x"e1",x"c0"),
   823 => (x"78",x"d4",x"48",x"d4"),
   824 => (x"48",x"ef",x"f1",x"c2"),
   825 => (x"50",x"bf",x"d4",x"ff"),
   826 => (x"ff",x"1e",x"4f",x"26"),
   827 => (x"e0",x"c0",x"48",x"d0"),
   828 => (x"1e",x"4f",x"26",x"78"),
   829 => (x"70",x"87",x"cc",x"ff"),
   830 => (x"c6",x"02",x"99",x"49"),
   831 => (x"a9",x"fb",x"c0",x"87"),
   832 => (x"71",x"87",x"f1",x"05"),
   833 => (x"0e",x"4f",x"26",x"48"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"4c",x"c0",x"4b",x"71"),
   836 => (x"70",x"87",x"f0",x"fe"),
   837 => (x"c0",x"02",x"99",x"49"),
   838 => (x"ec",x"c0",x"87",x"f9"),
   839 => (x"f2",x"c0",x"02",x"a9"),
   840 => (x"a9",x"fb",x"c0",x"87"),
   841 => (x"87",x"eb",x"c0",x"02"),
   842 => (x"ac",x"b7",x"66",x"cc"),
   843 => (x"d0",x"87",x"c7",x"03"),
   844 => (x"87",x"c2",x"02",x"66"),
   845 => (x"99",x"71",x"53",x"71"),
   846 => (x"c1",x"87",x"c2",x"02"),
   847 => (x"87",x"c3",x"fe",x"84"),
   848 => (x"02",x"99",x"49",x"70"),
   849 => (x"ec",x"c0",x"87",x"cd"),
   850 => (x"87",x"c7",x"02",x"a9"),
   851 => (x"05",x"a9",x"fb",x"c0"),
   852 => (x"d0",x"87",x"d5",x"ff"),
   853 => (x"87",x"c3",x"02",x"66"),
   854 => (x"c0",x"7b",x"97",x"c0"),
   855 => (x"c4",x"05",x"a9",x"ec"),
   856 => (x"c5",x"4a",x"74",x"87"),
   857 => (x"c0",x"4a",x"74",x"87"),
   858 => (x"48",x"72",x"8a",x"0a"),
   859 => (x"4d",x"26",x"87",x"c2"),
   860 => (x"4b",x"26",x"4c",x"26"),
   861 => (x"fd",x"1e",x"4f",x"26"),
   862 => (x"49",x"70",x"87",x"c9"),
   863 => (x"aa",x"f0",x"c0",x"4a"),
   864 => (x"c0",x"87",x"c9",x"04"),
   865 => (x"c3",x"01",x"aa",x"f9"),
   866 => (x"8a",x"f0",x"c0",x"87"),
   867 => (x"04",x"aa",x"c1",x"c1"),
   868 => (x"da",x"c1",x"87",x"c9"),
   869 => (x"87",x"c3",x"01",x"aa"),
   870 => (x"72",x"8a",x"f7",x"c0"),
   871 => (x"0e",x"4f",x"26",x"48"),
   872 => (x"0e",x"5c",x"5b",x"5e"),
   873 => (x"d4",x"ff",x"4a",x"71"),
   874 => (x"c0",x"49",x"72",x"4c"),
   875 => (x"4b",x"70",x"87",x"e9"),
   876 => (x"87",x"c2",x"02",x"9b"),
   877 => (x"d0",x"ff",x"8b",x"c1"),
   878 => (x"c1",x"78",x"c5",x"48"),
   879 => (x"49",x"73",x"7c",x"d5"),
   880 => (x"e7",x"c1",x"31",x"c6"),
   881 => (x"4a",x"bf",x"97",x"e2"),
   882 => (x"70",x"b0",x"71",x"48"),
   883 => (x"48",x"d0",x"ff",x"7c"),
   884 => (x"48",x"73",x"78",x"c4"),
   885 => (x"0e",x"87",x"d9",x"fe"),
   886 => (x"5d",x"5c",x"5b",x"5e"),
   887 => (x"71",x"86",x"f8",x"0e"),
   888 => (x"c0",x"7e",x"c0",x"4b"),
   889 => (x"bf",x"97",x"fe",x"fa"),
   890 => (x"05",x"a9",x"df",x"49"),
   891 => (x"c8",x"87",x"ee",x"c0"),
   892 => (x"69",x"97",x"49",x"a3"),
   893 => (x"a9",x"c3",x"c1",x"49"),
   894 => (x"c9",x"87",x"dd",x"05"),
   895 => (x"69",x"97",x"49",x"a3"),
   896 => (x"a9",x"c6",x"c1",x"49"),
   897 => (x"ca",x"87",x"d1",x"05"),
   898 => (x"69",x"97",x"49",x"a3"),
   899 => (x"a9",x"c7",x"c1",x"49"),
   900 => (x"c1",x"87",x"c5",x"05"),
   901 => (x"87",x"e1",x"c2",x"48"),
   902 => (x"dc",x"c2",x"48",x"c0"),
   903 => (x"87",x"ee",x"fa",x"87"),
   904 => (x"fa",x"c0",x"4c",x"c0"),
   905 => (x"49",x"bf",x"97",x"fe"),
   906 => (x"cf",x"04",x"a9",x"c0"),
   907 => (x"87",x"c3",x"fb",x"87"),
   908 => (x"fa",x"c0",x"84",x"c1"),
   909 => (x"49",x"bf",x"97",x"fe"),
   910 => (x"87",x"f1",x"06",x"ac"),
   911 => (x"97",x"fe",x"fa",x"c0"),
   912 => (x"87",x"cf",x"02",x"bf"),
   913 => (x"70",x"87",x"fc",x"f9"),
   914 => (x"c6",x"02",x"99",x"49"),
   915 => (x"a9",x"ec",x"c0",x"87"),
   916 => (x"c0",x"87",x"f1",x"05"),
   917 => (x"87",x"eb",x"f9",x"4c"),
   918 => (x"e6",x"f9",x"4d",x"70"),
   919 => (x"58",x"a6",x"c8",x"87"),
   920 => (x"70",x"87",x"e0",x"f9"),
   921 => (x"c8",x"84",x"c1",x"4a"),
   922 => (x"69",x"97",x"49",x"a3"),
   923 => (x"c7",x"02",x"ad",x"49"),
   924 => (x"ad",x"ff",x"c0",x"87"),
   925 => (x"87",x"e7",x"c0",x"05"),
   926 => (x"97",x"49",x"a3",x"c9"),
   927 => (x"66",x"c4",x"49",x"69"),
   928 => (x"87",x"c7",x"02",x"a9"),
   929 => (x"a8",x"ff",x"c0",x"48"),
   930 => (x"ca",x"87",x"d4",x"05"),
   931 => (x"69",x"97",x"49",x"a3"),
   932 => (x"c6",x"02",x"aa",x"49"),
   933 => (x"aa",x"ff",x"c0",x"87"),
   934 => (x"c1",x"87",x"c4",x"05"),
   935 => (x"c0",x"87",x"d0",x"7e"),
   936 => (x"c6",x"02",x"ad",x"ec"),
   937 => (x"ad",x"fb",x"c0",x"87"),
   938 => (x"c0",x"87",x"c4",x"05"),
   939 => (x"6e",x"7e",x"c1",x"4c"),
   940 => (x"87",x"e1",x"fe",x"02"),
   941 => (x"74",x"87",x"f3",x"f8"),
   942 => (x"fa",x"8e",x"f8",x"48"),
   943 => (x"0e",x"00",x"87",x"f0"),
   944 => (x"5d",x"5c",x"5b",x"5e"),
   945 => (x"71",x"86",x"f8",x"0e"),
   946 => (x"4b",x"d4",x"ff",x"4d"),
   947 => (x"f1",x"c2",x"1e",x"75"),
   948 => (x"ec",x"e4",x"49",x"f4"),
   949 => (x"70",x"86",x"c4",x"87"),
   950 => (x"cc",x"c4",x"02",x"98"),
   951 => (x"48",x"a6",x"c4",x"87"),
   952 => (x"bf",x"e4",x"e7",x"c1"),
   953 => (x"fa",x"49",x"75",x"78"),
   954 => (x"d0",x"ff",x"87",x"f5"),
   955 => (x"c1",x"78",x"c5",x"48"),
   956 => (x"4a",x"c0",x"7b",x"d6"),
   957 => (x"11",x"49",x"a2",x"75"),
   958 => (x"cb",x"82",x"c1",x"7b"),
   959 => (x"f3",x"04",x"aa",x"b7"),
   960 => (x"c3",x"4a",x"cc",x"87"),
   961 => (x"82",x"c1",x"7b",x"ff"),
   962 => (x"aa",x"b7",x"e0",x"c0"),
   963 => (x"ff",x"87",x"f4",x"04"),
   964 => (x"78",x"c4",x"48",x"d0"),
   965 => (x"c5",x"7b",x"ff",x"c3"),
   966 => (x"7b",x"d3",x"c1",x"78"),
   967 => (x"78",x"c4",x"7b",x"c1"),
   968 => (x"b7",x"c0",x"48",x"66"),
   969 => (x"f0",x"c2",x"06",x"a8"),
   970 => (x"fc",x"f1",x"c2",x"87"),
   971 => (x"66",x"c4",x"4c",x"bf"),
   972 => (x"c8",x"88",x"74",x"48"),
   973 => (x"9c",x"74",x"58",x"a6"),
   974 => (x"87",x"f9",x"c1",x"02"),
   975 => (x"7e",x"fe",x"e4",x"c2"),
   976 => (x"8c",x"4d",x"c0",x"c8"),
   977 => (x"03",x"ac",x"b7",x"c0"),
   978 => (x"c0",x"c8",x"87",x"c6"),
   979 => (x"4c",x"c0",x"4d",x"a4"),
   980 => (x"97",x"ef",x"f1",x"c2"),
   981 => (x"99",x"d0",x"49",x"bf"),
   982 => (x"c0",x"87",x"d1",x"02"),
   983 => (x"f4",x"f1",x"c2",x"1e"),
   984 => (x"87",x"d0",x"e7",x"49"),
   985 => (x"49",x"70",x"86",x"c4"),
   986 => (x"87",x"ee",x"c0",x"4a"),
   987 => (x"1e",x"fe",x"e4",x"c2"),
   988 => (x"49",x"f4",x"f1",x"c2"),
   989 => (x"c4",x"87",x"fd",x"e6"),
   990 => (x"4a",x"49",x"70",x"86"),
   991 => (x"c8",x"48",x"d0",x"ff"),
   992 => (x"d4",x"c1",x"78",x"c5"),
   993 => (x"bf",x"97",x"6e",x"7b"),
   994 => (x"c1",x"48",x"6e",x"7b"),
   995 => (x"c1",x"7e",x"70",x"80"),
   996 => (x"f0",x"ff",x"05",x"8d"),
   997 => (x"48",x"d0",x"ff",x"87"),
   998 => (x"9a",x"72",x"78",x"c4"),
   999 => (x"c0",x"87",x"c5",x"05"),
  1000 => (x"87",x"c7",x"c1",x"48"),
  1001 => (x"f1",x"c2",x"1e",x"c1"),
  1002 => (x"ed",x"e4",x"49",x"f4"),
  1003 => (x"74",x"86",x"c4",x"87"),
  1004 => (x"c7",x"fe",x"05",x"9c"),
  1005 => (x"48",x"66",x"c4",x"87"),
  1006 => (x"06",x"a8",x"b7",x"c0"),
  1007 => (x"f1",x"c2",x"87",x"d1"),
  1008 => (x"78",x"c0",x"48",x"f4"),
  1009 => (x"78",x"c0",x"80",x"d0"),
  1010 => (x"f2",x"c2",x"80",x"f4"),
  1011 => (x"c4",x"78",x"bf",x"c0"),
  1012 => (x"b7",x"c0",x"48",x"66"),
  1013 => (x"d0",x"fd",x"01",x"a8"),
  1014 => (x"48",x"d0",x"ff",x"87"),
  1015 => (x"d3",x"c1",x"78",x"c5"),
  1016 => (x"c4",x"7b",x"c0",x"7b"),
  1017 => (x"c2",x"48",x"c1",x"78"),
  1018 => (x"f8",x"48",x"c0",x"87"),
  1019 => (x"26",x"4d",x"26",x"8e"),
  1020 => (x"26",x"4b",x"26",x"4c"),
  1021 => (x"5b",x"5e",x"0e",x"4f"),
  1022 => (x"1e",x"0e",x"5d",x"5c"),
  1023 => (x"4c",x"c0",x"4b",x"71"),
  1024 => (x"c0",x"04",x"ab",x"4d"),
  1025 => (x"f7",x"c0",x"87",x"e8"),
  1026 => (x"9d",x"75",x"1e",x"d7"),
  1027 => (x"c0",x"87",x"c4",x"02"),
  1028 => (x"c1",x"87",x"c2",x"4a"),
  1029 => (x"ea",x"49",x"72",x"4a"),
  1030 => (x"86",x"c4",x"87",x"f0"),
  1031 => (x"84",x"c1",x"7e",x"70"),
  1032 => (x"87",x"c2",x"05",x"6e"),
  1033 => (x"85",x"c1",x"4c",x"73"),
  1034 => (x"ff",x"06",x"ac",x"73"),
  1035 => (x"48",x"6e",x"87",x"d8"),
  1036 => (x"87",x"f9",x"fe",x"26"),
  1037 => (x"5c",x"5b",x"5e",x"0e"),
  1038 => (x"cc",x"4b",x"71",x"0e"),
  1039 => (x"e8",x"c0",x"02",x"66"),
  1040 => (x"f0",x"c0",x"4c",x"87"),
  1041 => (x"e8",x"c0",x"02",x"8c"),
  1042 => (x"c1",x"4a",x"74",x"87"),
  1043 => (x"e0",x"c0",x"02",x"8a"),
  1044 => (x"dc",x"02",x"8a",x"87"),
  1045 => (x"d8",x"02",x"8a",x"87"),
  1046 => (x"8a",x"e0",x"c0",x"87"),
  1047 => (x"87",x"e5",x"c0",x"02"),
  1048 => (x"c0",x"02",x"8a",x"c1"),
  1049 => (x"ea",x"c0",x"87",x"e7"),
  1050 => (x"f9",x"49",x"73",x"87"),
  1051 => (x"e2",x"c0",x"87",x"d1"),
  1052 => (x"c0",x"1e",x"74",x"87"),
  1053 => (x"d8",x"db",x"c1",x"49"),
  1054 => (x"73",x"1e",x"74",x"87"),
  1055 => (x"d0",x"db",x"c1",x"49"),
  1056 => (x"ce",x"86",x"c8",x"87"),
  1057 => (x"c1",x"49",x"73",x"87"),
  1058 => (x"c6",x"87",x"e1",x"de"),
  1059 => (x"c1",x"49",x"73",x"87"),
  1060 => (x"fd",x"87",x"d1",x"df"),
  1061 => (x"5e",x"0e",x"87",x"d9"),
  1062 => (x"0e",x"5d",x"5c",x"5b"),
  1063 => (x"49",x"4c",x"71",x"1e"),
  1064 => (x"f2",x"c2",x"91",x"de"),
  1065 => (x"85",x"71",x"4d",x"dc"),
  1066 => (x"c1",x"02",x"6d",x"97"),
  1067 => (x"f2",x"c2",x"87",x"dd"),
  1068 => (x"74",x"4a",x"bf",x"c8"),
  1069 => (x"fc",x"49",x"72",x"82"),
  1070 => (x"7e",x"70",x"87",x"fb"),
  1071 => (x"f2",x"c0",x"02",x"6e"),
  1072 => (x"d0",x"f2",x"c2",x"87"),
  1073 => (x"cb",x"4a",x"6e",x"4b"),
  1074 => (x"db",x"ff",x"fe",x"49"),
  1075 => (x"cb",x"4b",x"74",x"87"),
  1076 => (x"d9",x"e8",x"c1",x"93"),
  1077 => (x"c1",x"83",x"c4",x"83"),
  1078 => (x"74",x"7b",x"cf",x"c4"),
  1079 => (x"c9",x"c5",x"c1",x"49"),
  1080 => (x"c1",x"7b",x"75",x"87"),
  1081 => (x"bf",x"97",x"e3",x"e7"),
  1082 => (x"f2",x"c2",x"1e",x"49"),
  1083 => (x"c3",x"fd",x"49",x"d0"),
  1084 => (x"74",x"86",x"c4",x"87"),
  1085 => (x"f1",x"c4",x"c1",x"49"),
  1086 => (x"c1",x"49",x"c0",x"87"),
  1087 => (x"c2",x"87",x"d0",x"c6"),
  1088 => (x"c0",x"48",x"f0",x"f1"),
  1089 => (x"c0",x"49",x"c1",x"78"),
  1090 => (x"26",x"87",x"cf",x"e0"),
  1091 => (x"4c",x"87",x"de",x"fb"),
  1092 => (x"69",x"64",x"61",x"6f"),
  1093 => (x"2e",x"2e",x"67",x"6e"),
  1094 => (x"5e",x"0e",x"00",x"2e"),
  1095 => (x"71",x"0e",x"5c",x"5b"),
  1096 => (x"f2",x"c2",x"4a",x"4b"),
  1097 => (x"72",x"82",x"bf",x"c8"),
  1098 => (x"87",x"c9",x"fb",x"49"),
  1099 => (x"02",x"9c",x"4c",x"70"),
  1100 => (x"e5",x"49",x"87",x"c4"),
  1101 => (x"f2",x"c2",x"87",x"dc"),
  1102 => (x"78",x"c0",x"48",x"c8"),
  1103 => (x"d9",x"df",x"49",x"c1"),
  1104 => (x"87",x"eb",x"fa",x"87"),
  1105 => (x"5c",x"5b",x"5e",x"0e"),
  1106 => (x"86",x"f4",x"0e",x"5d"),
  1107 => (x"4d",x"fe",x"e4",x"c2"),
  1108 => (x"a6",x"c4",x"4c",x"c0"),
  1109 => (x"c2",x"78",x"c0",x"48"),
  1110 => (x"49",x"bf",x"c8",x"f2"),
  1111 => (x"c1",x"06",x"a9",x"c0"),
  1112 => (x"e4",x"c2",x"87",x"c1"),
  1113 => (x"02",x"98",x"48",x"fe"),
  1114 => (x"c0",x"87",x"f8",x"c0"),
  1115 => (x"c8",x"1e",x"d7",x"f7"),
  1116 => (x"87",x"c7",x"02",x"66"),
  1117 => (x"c0",x"48",x"a6",x"c4"),
  1118 => (x"c4",x"87",x"c5",x"78"),
  1119 => (x"78",x"c1",x"48",x"a6"),
  1120 => (x"e5",x"49",x"66",x"c4"),
  1121 => (x"86",x"c4",x"87",x"c4"),
  1122 => (x"84",x"c1",x"4d",x"70"),
  1123 => (x"c1",x"48",x"66",x"c4"),
  1124 => (x"58",x"a6",x"c8",x"80"),
  1125 => (x"bf",x"c8",x"f2",x"c2"),
  1126 => (x"c6",x"03",x"ac",x"49"),
  1127 => (x"05",x"9d",x"75",x"87"),
  1128 => (x"c0",x"87",x"c8",x"ff"),
  1129 => (x"02",x"9d",x"75",x"4c"),
  1130 => (x"c0",x"87",x"e0",x"c3"),
  1131 => (x"c8",x"1e",x"d7",x"f7"),
  1132 => (x"87",x"c7",x"02",x"66"),
  1133 => (x"c0",x"48",x"a6",x"cc"),
  1134 => (x"cc",x"87",x"c5",x"78"),
  1135 => (x"78",x"c1",x"48",x"a6"),
  1136 => (x"e4",x"49",x"66",x"cc"),
  1137 => (x"86",x"c4",x"87",x"c4"),
  1138 => (x"02",x"6e",x"7e",x"70"),
  1139 => (x"6e",x"87",x"e9",x"c2"),
  1140 => (x"97",x"81",x"cb",x"49"),
  1141 => (x"99",x"d0",x"49",x"69"),
  1142 => (x"87",x"d6",x"c1",x"02"),
  1143 => (x"4a",x"da",x"c4",x"c1"),
  1144 => (x"91",x"cb",x"49",x"74"),
  1145 => (x"81",x"d9",x"e8",x"c1"),
  1146 => (x"81",x"c8",x"79",x"72"),
  1147 => (x"74",x"51",x"ff",x"c3"),
  1148 => (x"c2",x"91",x"de",x"49"),
  1149 => (x"71",x"4d",x"dc",x"f2"),
  1150 => (x"97",x"c1",x"c2",x"85"),
  1151 => (x"49",x"a5",x"c1",x"7d"),
  1152 => (x"c2",x"51",x"e0",x"c0"),
  1153 => (x"bf",x"97",x"ce",x"ed"),
  1154 => (x"c1",x"87",x"d2",x"02"),
  1155 => (x"4b",x"a5",x"c2",x"84"),
  1156 => (x"4a",x"ce",x"ed",x"c2"),
  1157 => (x"fa",x"fe",x"49",x"db"),
  1158 => (x"db",x"c1",x"87",x"ce"),
  1159 => (x"49",x"a5",x"cd",x"87"),
  1160 => (x"84",x"c1",x"51",x"c0"),
  1161 => (x"6e",x"4b",x"a5",x"c2"),
  1162 => (x"fe",x"49",x"cb",x"4a"),
  1163 => (x"c1",x"87",x"f9",x"f9"),
  1164 => (x"c2",x"c1",x"87",x"c6"),
  1165 => (x"49",x"74",x"4a",x"d6"),
  1166 => (x"e8",x"c1",x"91",x"cb"),
  1167 => (x"79",x"72",x"81",x"d9"),
  1168 => (x"97",x"ce",x"ed",x"c2"),
  1169 => (x"87",x"d8",x"02",x"bf"),
  1170 => (x"91",x"de",x"49",x"74"),
  1171 => (x"f2",x"c2",x"84",x"c1"),
  1172 => (x"83",x"71",x"4b",x"dc"),
  1173 => (x"4a",x"ce",x"ed",x"c2"),
  1174 => (x"f9",x"fe",x"49",x"dd"),
  1175 => (x"87",x"d8",x"87",x"ca"),
  1176 => (x"93",x"de",x"4b",x"74"),
  1177 => (x"83",x"dc",x"f2",x"c2"),
  1178 => (x"c0",x"49",x"a3",x"cb"),
  1179 => (x"73",x"84",x"c1",x"51"),
  1180 => (x"49",x"cb",x"4a",x"6e"),
  1181 => (x"87",x"f0",x"f8",x"fe"),
  1182 => (x"c1",x"48",x"66",x"c4"),
  1183 => (x"58",x"a6",x"c8",x"80"),
  1184 => (x"c0",x"03",x"ac",x"c7"),
  1185 => (x"05",x"6e",x"87",x"c5"),
  1186 => (x"74",x"87",x"e0",x"fc"),
  1187 => (x"f5",x"8e",x"f4",x"48"),
  1188 => (x"73",x"1e",x"87",x"db"),
  1189 => (x"49",x"4b",x"71",x"1e"),
  1190 => (x"e8",x"c1",x"91",x"cb"),
  1191 => (x"a1",x"c8",x"81",x"d9"),
  1192 => (x"e2",x"e7",x"c1",x"4a"),
  1193 => (x"c9",x"50",x"12",x"48"),
  1194 => (x"fa",x"c0",x"4a",x"a1"),
  1195 => (x"50",x"12",x"48",x"fe"),
  1196 => (x"e7",x"c1",x"81",x"ca"),
  1197 => (x"50",x"11",x"48",x"e3"),
  1198 => (x"97",x"e3",x"e7",x"c1"),
  1199 => (x"c0",x"1e",x"49",x"bf"),
  1200 => (x"87",x"f0",x"f5",x"49"),
  1201 => (x"48",x"f0",x"f1",x"c2"),
  1202 => (x"49",x"c1",x"78",x"de"),
  1203 => (x"26",x"87",x"cb",x"d9"),
  1204 => (x"1e",x"87",x"de",x"f4"),
  1205 => (x"cb",x"49",x"4a",x"71"),
  1206 => (x"d9",x"e8",x"c1",x"91"),
  1207 => (x"11",x"81",x"c8",x"81"),
  1208 => (x"f4",x"f1",x"c2",x"48"),
  1209 => (x"c8",x"f2",x"c2",x"58"),
  1210 => (x"c1",x"78",x"c0",x"48"),
  1211 => (x"87",x"ea",x"d8",x"49"),
  1212 => (x"c0",x"1e",x"4f",x"26"),
  1213 => (x"d6",x"fe",x"c0",x"49"),
  1214 => (x"1e",x"4f",x"26",x"87"),
  1215 => (x"d2",x"02",x"99",x"71"),
  1216 => (x"ee",x"e9",x"c1",x"87"),
  1217 => (x"f7",x"50",x"c0",x"48"),
  1218 => (x"d3",x"cb",x"c1",x"80"),
  1219 => (x"c7",x"e8",x"c1",x"40"),
  1220 => (x"c1",x"87",x"ce",x"78"),
  1221 => (x"c1",x"48",x"ea",x"e9"),
  1222 => (x"fc",x"78",x"e8",x"e7"),
  1223 => (x"f2",x"cb",x"c1",x"80"),
  1224 => (x"0e",x"4f",x"26",x"78"),
  1225 => (x"0e",x"5c",x"5b",x"5e"),
  1226 => (x"cb",x"4a",x"4c",x"71"),
  1227 => (x"d9",x"e8",x"c1",x"92"),
  1228 => (x"49",x"a2",x"c8",x"82"),
  1229 => (x"97",x"4b",x"a2",x"c9"),
  1230 => (x"97",x"1e",x"4b",x"6b"),
  1231 => (x"ca",x"1e",x"49",x"69"),
  1232 => (x"c0",x"49",x"12",x"82"),
  1233 => (x"c0",x"87",x"d1",x"e9"),
  1234 => (x"87",x"ce",x"d7",x"49"),
  1235 => (x"fb",x"c0",x"49",x"74"),
  1236 => (x"8e",x"f8",x"87",x"d8"),
  1237 => (x"1e",x"87",x"d8",x"f2"),
  1238 => (x"4b",x"71",x"1e",x"73"),
  1239 => (x"87",x"c3",x"ff",x"49"),
  1240 => (x"fe",x"fe",x"49",x"73"),
  1241 => (x"c0",x"49",x"c0",x"87"),
  1242 => (x"f2",x"87",x"e4",x"fc"),
  1243 => (x"73",x"1e",x"87",x"c3"),
  1244 => (x"c6",x"4b",x"71",x"1e"),
  1245 => (x"dc",x"02",x"4a",x"a3"),
  1246 => (x"02",x"8a",x"c1",x"87"),
  1247 => (x"8a",x"87",x"e4",x"c0"),
  1248 => (x"87",x"e8",x"c1",x"02"),
  1249 => (x"ca",x"c1",x"02",x"8a"),
  1250 => (x"c0",x"02",x"8a",x"87"),
  1251 => (x"02",x"8a",x"87",x"ef"),
  1252 => (x"e9",x"c1",x"87",x"d9"),
  1253 => (x"f0",x"f1",x"c2",x"87"),
  1254 => (x"c1",x"78",x"df",x"48"),
  1255 => (x"87",x"fa",x"d5",x"49"),
  1256 => (x"c7",x"87",x"e6",x"c1"),
  1257 => (x"87",x"eb",x"fc",x"49"),
  1258 => (x"c2",x"87",x"de",x"c1"),
  1259 => (x"02",x"bf",x"c8",x"f2"),
  1260 => (x"48",x"87",x"cb",x"c1"),
  1261 => (x"f2",x"c2",x"88",x"c1"),
  1262 => (x"c1",x"c1",x"58",x"cc"),
  1263 => (x"cc",x"f2",x"c2",x"87"),
  1264 => (x"f9",x"c0",x"02",x"bf"),
  1265 => (x"c8",x"f2",x"c2",x"87"),
  1266 => (x"80",x"c1",x"48",x"bf"),
  1267 => (x"58",x"cc",x"f2",x"c2"),
  1268 => (x"c2",x"87",x"eb",x"c0"),
  1269 => (x"49",x"bf",x"c8",x"f2"),
  1270 => (x"f2",x"c2",x"89",x"c6"),
  1271 => (x"b7",x"c0",x"59",x"cc"),
  1272 => (x"87",x"da",x"03",x"a9"),
  1273 => (x"48",x"c8",x"f2",x"c2"),
  1274 => (x"87",x"d2",x"78",x"c0"),
  1275 => (x"bf",x"cc",x"f2",x"c2"),
  1276 => (x"c2",x"87",x"cb",x"02"),
  1277 => (x"48",x"bf",x"c8",x"f2"),
  1278 => (x"f2",x"c2",x"80",x"c6"),
  1279 => (x"49",x"c0",x"58",x"cc"),
  1280 => (x"73",x"87",x"d7",x"d4"),
  1281 => (x"e1",x"f8",x"c0",x"49"),
  1282 => (x"87",x"e5",x"ef",x"87"),
  1283 => (x"5c",x"5b",x"5e",x"0e"),
  1284 => (x"d0",x"ff",x"0e",x"5d"),
  1285 => (x"59",x"a6",x"dc",x"86"),
  1286 => (x"c0",x"48",x"a6",x"c8"),
  1287 => (x"c1",x"80",x"c4",x"78"),
  1288 => (x"c4",x"78",x"66",x"c4"),
  1289 => (x"c4",x"78",x"c1",x"80"),
  1290 => (x"c2",x"78",x"c1",x"80"),
  1291 => (x"c1",x"48",x"cc",x"f2"),
  1292 => (x"f0",x"f1",x"c2",x"78"),
  1293 => (x"48",x"6e",x"7e",x"bf"),
  1294 => (x"cb",x"05",x"a8",x"de"),
  1295 => (x"87",x"c4",x"f4",x"87"),
  1296 => (x"a6",x"cc",x"49",x"70"),
  1297 => (x"87",x"f1",x"d1",x"59"),
  1298 => (x"a8",x"df",x"48",x"6e"),
  1299 => (x"87",x"ee",x"c1",x"05"),
  1300 => (x"49",x"66",x"c0",x"c1"),
  1301 => (x"7e",x"69",x"81",x"c4"),
  1302 => (x"48",x"ee",x"e3",x"c1"),
  1303 => (x"a1",x"d0",x"49",x"6e"),
  1304 => (x"71",x"41",x"20",x"4a"),
  1305 => (x"87",x"f9",x"05",x"aa"),
  1306 => (x"4a",x"d2",x"ca",x"c1"),
  1307 => (x"0a",x"66",x"c0",x"c1"),
  1308 => (x"c0",x"c1",x"0a",x"7a"),
  1309 => (x"81",x"c9",x"49",x"66"),
  1310 => (x"c0",x"c1",x"51",x"df"),
  1311 => (x"81",x"ca",x"49",x"66"),
  1312 => (x"c1",x"51",x"d3",x"c1"),
  1313 => (x"cb",x"49",x"66",x"c0"),
  1314 => (x"4b",x"a1",x"c4",x"81"),
  1315 => (x"6b",x"48",x"a6",x"c4"),
  1316 => (x"72",x"1e",x"71",x"78"),
  1317 => (x"fe",x"e3",x"c1",x"1e"),
  1318 => (x"49",x"66",x"cc",x"48"),
  1319 => (x"20",x"4a",x"a1",x"d0"),
  1320 => (x"05",x"aa",x"71",x"41"),
  1321 => (x"4a",x"26",x"87",x"f9"),
  1322 => (x"79",x"72",x"49",x"26"),
  1323 => (x"df",x"4a",x"a1",x"c9"),
  1324 => (x"c1",x"81",x"ca",x"52"),
  1325 => (x"a6",x"c8",x"51",x"d4"),
  1326 => (x"cf",x"78",x"c2",x"48"),
  1327 => (x"cd",x"e0",x"87",x"fb"),
  1328 => (x"87",x"ef",x"e0",x"87"),
  1329 => (x"87",x"fb",x"df",x"ff"),
  1330 => (x"fb",x"c0",x"4c",x"70"),
  1331 => (x"fd",x"c1",x"02",x"ac"),
  1332 => (x"05",x"66",x"d8",x"87"),
  1333 => (x"c1",x"87",x"ee",x"c1"),
  1334 => (x"c4",x"4a",x"66",x"c0"),
  1335 => (x"72",x"7e",x"6a",x"82"),
  1336 => (x"ce",x"e4",x"c1",x"1e"),
  1337 => (x"49",x"66",x"c4",x"48"),
  1338 => (x"20",x"4a",x"a1",x"c8"),
  1339 => (x"05",x"aa",x"71",x"41"),
  1340 => (x"51",x"10",x"87",x"f9"),
  1341 => (x"c0",x"c1",x"4a",x"26"),
  1342 => (x"ca",x"c1",x"48",x"66"),
  1343 => (x"49",x"6a",x"78",x"d2"),
  1344 => (x"51",x"74",x"81",x"c7"),
  1345 => (x"49",x"66",x"c0",x"c1"),
  1346 => (x"51",x"c1",x"81",x"c8"),
  1347 => (x"49",x"66",x"c0",x"c1"),
  1348 => (x"51",x"c0",x"81",x"c9"),
  1349 => (x"49",x"66",x"c0",x"c1"),
  1350 => (x"51",x"c0",x"81",x"ca"),
  1351 => (x"1e",x"d8",x"1e",x"c1"),
  1352 => (x"81",x"c8",x"49",x"6a"),
  1353 => (x"87",x"df",x"df",x"ff"),
  1354 => (x"c4",x"c1",x"86",x"c8"),
  1355 => (x"a8",x"c0",x"48",x"66"),
  1356 => (x"c8",x"87",x"c7",x"01"),
  1357 => (x"78",x"c1",x"48",x"a6"),
  1358 => (x"c4",x"c1",x"87",x"cf"),
  1359 => (x"88",x"c1",x"48",x"66"),
  1360 => (x"c4",x"58",x"a6",x"d0"),
  1361 => (x"ea",x"de",x"ff",x"87"),
  1362 => (x"48",x"a6",x"d0",x"87"),
  1363 => (x"9c",x"74",x"78",x"c2"),
  1364 => (x"87",x"e1",x"cd",x"02"),
  1365 => (x"c1",x"48",x"66",x"c8"),
  1366 => (x"03",x"a8",x"66",x"c8"),
  1367 => (x"dc",x"87",x"d6",x"cd"),
  1368 => (x"78",x"c0",x"48",x"a6"),
  1369 => (x"78",x"c0",x"80",x"e8"),
  1370 => (x"87",x"d7",x"dd",x"ff"),
  1371 => (x"d0",x"c1",x"4c",x"70"),
  1372 => (x"db",x"c2",x"05",x"ac"),
  1373 => (x"7e",x"66",x"c4",x"87"),
  1374 => (x"87",x"fa",x"df",x"ff"),
  1375 => (x"a6",x"c8",x"49",x"70"),
  1376 => (x"fe",x"dc",x"ff",x"59"),
  1377 => (x"c0",x"4c",x"70",x"87"),
  1378 => (x"c1",x"05",x"ac",x"ec"),
  1379 => (x"66",x"c8",x"87",x"ed"),
  1380 => (x"c1",x"91",x"cb",x"49"),
  1381 => (x"c4",x"81",x"66",x"c0"),
  1382 => (x"4d",x"6a",x"4a",x"a1"),
  1383 => (x"c4",x"4a",x"a1",x"c8"),
  1384 => (x"cb",x"c1",x"52",x"66"),
  1385 => (x"dc",x"ff",x"79",x"d3"),
  1386 => (x"4c",x"70",x"87",x"d9"),
  1387 => (x"87",x"d9",x"02",x"9c"),
  1388 => (x"02",x"ac",x"fb",x"c0"),
  1389 => (x"55",x"74",x"87",x"d3"),
  1390 => (x"87",x"c7",x"dc",x"ff"),
  1391 => (x"02",x"9c",x"4c",x"70"),
  1392 => (x"fb",x"c0",x"87",x"c7"),
  1393 => (x"ed",x"ff",x"05",x"ac"),
  1394 => (x"55",x"e0",x"c0",x"87"),
  1395 => (x"c0",x"55",x"c1",x"c2"),
  1396 => (x"66",x"d8",x"7d",x"97"),
  1397 => (x"05",x"a9",x"6e",x"49"),
  1398 => (x"66",x"c8",x"87",x"db"),
  1399 => (x"a8",x"66",x"cc",x"48"),
  1400 => (x"c8",x"87",x"ca",x"04"),
  1401 => (x"80",x"c1",x"48",x"66"),
  1402 => (x"c8",x"58",x"a6",x"cc"),
  1403 => (x"48",x"66",x"cc",x"87"),
  1404 => (x"a6",x"d0",x"88",x"c1"),
  1405 => (x"ca",x"db",x"ff",x"58"),
  1406 => (x"c1",x"4c",x"70",x"87"),
  1407 => (x"c8",x"05",x"ac",x"d0"),
  1408 => (x"48",x"66",x"d4",x"87"),
  1409 => (x"a6",x"d8",x"80",x"c1"),
  1410 => (x"ac",x"d0",x"c1",x"58"),
  1411 => (x"87",x"e5",x"fd",x"02"),
  1412 => (x"48",x"a6",x"e0",x"c0"),
  1413 => (x"c4",x"78",x"66",x"d8"),
  1414 => (x"e0",x"c0",x"48",x"66"),
  1415 => (x"c9",x"05",x"a8",x"66"),
  1416 => (x"e4",x"c0",x"87",x"e5"),
  1417 => (x"78",x"c0",x"48",x"a6"),
  1418 => (x"78",x"c0",x"80",x"c4"),
  1419 => (x"fb",x"c0",x"48",x"74"),
  1420 => (x"6e",x"7e",x"70",x"88"),
  1421 => (x"87",x"e8",x"c8",x"02"),
  1422 => (x"88",x"cb",x"48",x"6e"),
  1423 => (x"02",x"6e",x"7e",x"70"),
  1424 => (x"6e",x"87",x"ce",x"c1"),
  1425 => (x"70",x"88",x"c9",x"48"),
  1426 => (x"c3",x"02",x"6e",x"7e"),
  1427 => (x"48",x"6e",x"87",x"ea"),
  1428 => (x"7e",x"70",x"88",x"c4"),
  1429 => (x"87",x"ce",x"02",x"6e"),
  1430 => (x"88",x"c1",x"48",x"6e"),
  1431 => (x"02",x"6e",x"7e",x"70"),
  1432 => (x"c7",x"87",x"d5",x"c3"),
  1433 => (x"a6",x"dc",x"87",x"f4"),
  1434 => (x"78",x"f0",x"c0",x"48"),
  1435 => (x"87",x"d3",x"d9",x"ff"),
  1436 => (x"ec",x"c0",x"4c",x"70"),
  1437 => (x"c4",x"c0",x"02",x"ac"),
  1438 => (x"a6",x"e0",x"c0",x"87"),
  1439 => (x"ac",x"ec",x"c0",x"5c"),
  1440 => (x"87",x"cd",x"c0",x"02"),
  1441 => (x"87",x"fb",x"d8",x"ff"),
  1442 => (x"ec",x"c0",x"4c",x"70"),
  1443 => (x"f3",x"ff",x"05",x"ac"),
  1444 => (x"ac",x"ec",x"c0",x"87"),
  1445 => (x"87",x"c4",x"c0",x"02"),
  1446 => (x"87",x"e7",x"d8",x"ff"),
  1447 => (x"1e",x"ca",x"1e",x"c0"),
  1448 => (x"cb",x"49",x"66",x"d0"),
  1449 => (x"66",x"c8",x"c1",x"91"),
  1450 => (x"cc",x"80",x"71",x"48"),
  1451 => (x"66",x"c8",x"58",x"a6"),
  1452 => (x"d0",x"80",x"c4",x"48"),
  1453 => (x"66",x"cc",x"58",x"a6"),
  1454 => (x"d9",x"ff",x"49",x"bf"),
  1455 => (x"1e",x"c1",x"87",x"c9"),
  1456 => (x"66",x"d4",x"1e",x"de"),
  1457 => (x"d8",x"ff",x"49",x"bf"),
  1458 => (x"86",x"d0",x"87",x"fd"),
  1459 => (x"09",x"c0",x"49",x"70"),
  1460 => (x"a6",x"ec",x"c0",x"89"),
  1461 => (x"66",x"e8",x"c0",x"59"),
  1462 => (x"06",x"a8",x"c0",x"48"),
  1463 => (x"c0",x"87",x"ee",x"c0"),
  1464 => (x"dd",x"48",x"66",x"e8"),
  1465 => (x"e4",x"c0",x"03",x"a8"),
  1466 => (x"bf",x"66",x"c4",x"87"),
  1467 => (x"66",x"e8",x"c0",x"49"),
  1468 => (x"51",x"e0",x"c0",x"81"),
  1469 => (x"49",x"66",x"e8",x"c0"),
  1470 => (x"66",x"c4",x"81",x"c1"),
  1471 => (x"c1",x"c2",x"81",x"bf"),
  1472 => (x"66",x"e8",x"c0",x"51"),
  1473 => (x"c4",x"81",x"c2",x"49"),
  1474 => (x"c0",x"81",x"bf",x"66"),
  1475 => (x"c1",x"48",x"6e",x"51"),
  1476 => (x"6e",x"78",x"d2",x"ca"),
  1477 => (x"d0",x"81",x"c8",x"49"),
  1478 => (x"49",x"6e",x"51",x"66"),
  1479 => (x"66",x"d4",x"81",x"c9"),
  1480 => (x"ca",x"49",x"6e",x"51"),
  1481 => (x"51",x"66",x"dc",x"81"),
  1482 => (x"c1",x"48",x"66",x"d0"),
  1483 => (x"58",x"a6",x"d4",x"80"),
  1484 => (x"c1",x"80",x"d8",x"48"),
  1485 => (x"87",x"e8",x"c4",x"78"),
  1486 => (x"87",x"fa",x"d8",x"ff"),
  1487 => (x"ec",x"c0",x"49",x"70"),
  1488 => (x"d8",x"ff",x"59",x"a6"),
  1489 => (x"49",x"70",x"87",x"f0"),
  1490 => (x"59",x"a6",x"e0",x"c0"),
  1491 => (x"c0",x"48",x"66",x"dc"),
  1492 => (x"c0",x"05",x"a8",x"ec"),
  1493 => (x"a6",x"dc",x"87",x"ca"),
  1494 => (x"66",x"e8",x"c0",x"48"),
  1495 => (x"87",x"c4",x"c0",x"78"),
  1496 => (x"87",x"df",x"d5",x"ff"),
  1497 => (x"cb",x"49",x"66",x"c8"),
  1498 => (x"66",x"c0",x"c1",x"91"),
  1499 => (x"70",x"80",x"71",x"48"),
  1500 => (x"c8",x"4a",x"6e",x"7e"),
  1501 => (x"ca",x"49",x"6e",x"82"),
  1502 => (x"66",x"e8",x"c0",x"81"),
  1503 => (x"49",x"66",x"dc",x"51"),
  1504 => (x"e8",x"c0",x"81",x"c1"),
  1505 => (x"48",x"c1",x"89",x"66"),
  1506 => (x"49",x"70",x"30",x"71"),
  1507 => (x"97",x"71",x"89",x"c1"),
  1508 => (x"f8",x"f5",x"c2",x"7a"),
  1509 => (x"e8",x"c0",x"49",x"bf"),
  1510 => (x"6a",x"97",x"29",x"66"),
  1511 => (x"98",x"71",x"48",x"4a"),
  1512 => (x"58",x"a6",x"f0",x"c0"),
  1513 => (x"81",x"c4",x"49",x"6e"),
  1514 => (x"e0",x"c0",x"4d",x"69"),
  1515 => (x"66",x"c4",x"48",x"66"),
  1516 => (x"c8",x"c0",x"02",x"a8"),
  1517 => (x"48",x"a6",x"c4",x"87"),
  1518 => (x"c5",x"c0",x"78",x"c0"),
  1519 => (x"48",x"a6",x"c4",x"87"),
  1520 => (x"66",x"c4",x"78",x"c1"),
  1521 => (x"1e",x"e0",x"c0",x"1e"),
  1522 => (x"d4",x"ff",x"49",x"75"),
  1523 => (x"86",x"c8",x"87",x"f9"),
  1524 => (x"b7",x"c0",x"4c",x"70"),
  1525 => (x"d4",x"c1",x"06",x"ac"),
  1526 => (x"c0",x"85",x"74",x"87"),
  1527 => (x"89",x"74",x"49",x"e0"),
  1528 => (x"e4",x"c1",x"4b",x"75"),
  1529 => (x"fe",x"71",x"4a",x"d7"),
  1530 => (x"c2",x"87",x"fd",x"e2"),
  1531 => (x"66",x"e4",x"c0",x"85"),
  1532 => (x"c0",x"80",x"c1",x"48"),
  1533 => (x"c0",x"58",x"a6",x"e8"),
  1534 => (x"c1",x"49",x"66",x"ec"),
  1535 => (x"02",x"a9",x"70",x"81"),
  1536 => (x"c4",x"87",x"c8",x"c0"),
  1537 => (x"78",x"c0",x"48",x"a6"),
  1538 => (x"c4",x"87",x"c5",x"c0"),
  1539 => (x"78",x"c1",x"48",x"a6"),
  1540 => (x"c2",x"1e",x"66",x"c4"),
  1541 => (x"e0",x"c0",x"49",x"a4"),
  1542 => (x"70",x"88",x"71",x"48"),
  1543 => (x"49",x"75",x"1e",x"49"),
  1544 => (x"87",x"e3",x"d3",x"ff"),
  1545 => (x"b7",x"c0",x"86",x"c8"),
  1546 => (x"c0",x"ff",x"01",x"a8"),
  1547 => (x"66",x"e4",x"c0",x"87"),
  1548 => (x"87",x"d1",x"c0",x"02"),
  1549 => (x"81",x"c9",x"49",x"6e"),
  1550 => (x"51",x"66",x"e4",x"c0"),
  1551 => (x"cc",x"c1",x"48",x"6e"),
  1552 => (x"cc",x"c0",x"78",x"e3"),
  1553 => (x"c9",x"49",x"6e",x"87"),
  1554 => (x"6e",x"51",x"c2",x"81"),
  1555 => (x"d7",x"cd",x"c1",x"48"),
  1556 => (x"a6",x"e8",x"c0",x"78"),
  1557 => (x"c0",x"78",x"c1",x"48"),
  1558 => (x"d2",x"ff",x"87",x"c6"),
  1559 => (x"4c",x"70",x"87",x"d5"),
  1560 => (x"02",x"66",x"e8",x"c0"),
  1561 => (x"c8",x"87",x"f5",x"c0"),
  1562 => (x"66",x"cc",x"48",x"66"),
  1563 => (x"cb",x"c0",x"04",x"a8"),
  1564 => (x"48",x"66",x"c8",x"87"),
  1565 => (x"a6",x"cc",x"80",x"c1"),
  1566 => (x"87",x"e0",x"c0",x"58"),
  1567 => (x"c1",x"48",x"66",x"cc"),
  1568 => (x"58",x"a6",x"d0",x"88"),
  1569 => (x"c1",x"87",x"d5",x"c0"),
  1570 => (x"c0",x"05",x"ac",x"c6"),
  1571 => (x"66",x"d0",x"87",x"c8"),
  1572 => (x"d4",x"80",x"c1",x"48"),
  1573 => (x"d1",x"ff",x"58",x"a6"),
  1574 => (x"4c",x"70",x"87",x"d9"),
  1575 => (x"c1",x"48",x"66",x"d4"),
  1576 => (x"58",x"a6",x"d8",x"80"),
  1577 => (x"c0",x"02",x"9c",x"74"),
  1578 => (x"66",x"c8",x"87",x"cb"),
  1579 => (x"66",x"c8",x"c1",x"48"),
  1580 => (x"ea",x"f2",x"04",x"a8"),
  1581 => (x"f1",x"d0",x"ff",x"87"),
  1582 => (x"48",x"66",x"c8",x"87"),
  1583 => (x"c0",x"03",x"a8",x"c7"),
  1584 => (x"f2",x"c2",x"87",x"e5"),
  1585 => (x"78",x"c0",x"48",x"cc"),
  1586 => (x"cb",x"49",x"66",x"c8"),
  1587 => (x"66",x"c0",x"c1",x"91"),
  1588 => (x"4a",x"a1",x"c4",x"81"),
  1589 => (x"52",x"c0",x"4a",x"6a"),
  1590 => (x"48",x"66",x"c8",x"79"),
  1591 => (x"a6",x"cc",x"80",x"c1"),
  1592 => (x"04",x"a8",x"c7",x"58"),
  1593 => (x"ff",x"87",x"db",x"ff"),
  1594 => (x"db",x"ff",x"8e",x"d0"),
  1595 => (x"6f",x"4c",x"87",x"ff"),
  1596 => (x"53",x"20",x"64",x"61"),
  1597 => (x"69",x"74",x"74",x"65"),
  1598 => (x"20",x"73",x"67",x"6e"),
  1599 => (x"61",x"53",x"00",x"81"),
  1600 => (x"53",x"20",x"65",x"76"),
  1601 => (x"69",x"74",x"74",x"65"),
  1602 => (x"20",x"73",x"67",x"6e"),
  1603 => (x"6f",x"4c",x"00",x"81"),
  1604 => (x"2a",x"20",x"64",x"61"),
  1605 => (x"3a",x"00",x"20",x"2e"),
  1606 => (x"73",x"1e",x"00",x"20"),
  1607 => (x"9b",x"4b",x"71",x"1e"),
  1608 => (x"c2",x"87",x"c6",x"02"),
  1609 => (x"c0",x"48",x"c8",x"f2"),
  1610 => (x"c2",x"1e",x"c7",x"78"),
  1611 => (x"49",x"bf",x"c8",x"f2"),
  1612 => (x"d9",x"e8",x"c1",x"1e"),
  1613 => (x"f0",x"f1",x"c2",x"1e"),
  1614 => (x"cf",x"eb",x"49",x"bf"),
  1615 => (x"c2",x"86",x"cc",x"87"),
  1616 => (x"49",x"bf",x"f0",x"f1"),
  1617 => (x"73",x"87",x"f4",x"e6"),
  1618 => (x"87",x"c8",x"02",x"9b"),
  1619 => (x"49",x"d9",x"e8",x"c1"),
  1620 => (x"87",x"e8",x"e4",x"c0"),
  1621 => (x"87",x"d9",x"da",x"ff"),
  1622 => (x"87",x"f7",x"c7",x"1e"),
  1623 => (x"f9",x"fe",x"49",x"c1"),
  1624 => (x"eb",x"e5",x"fe",x"87"),
  1625 => (x"02",x"98",x"70",x"87"),
  1626 => (x"ee",x"fe",x"87",x"cd"),
  1627 => (x"98",x"70",x"87",x"e6"),
  1628 => (x"c1",x"87",x"c4",x"02"),
  1629 => (x"c0",x"87",x"c2",x"4a"),
  1630 => (x"05",x"9a",x"72",x"4a"),
  1631 => (x"1e",x"c0",x"87",x"ce"),
  1632 => (x"49",x"e9",x"e6",x"c1"),
  1633 => (x"87",x"c3",x"f0",x"c0"),
  1634 => (x"87",x"fe",x"86",x"c4"),
  1635 => (x"e6",x"c1",x"1e",x"c0"),
  1636 => (x"ef",x"c0",x"49",x"f4"),
  1637 => (x"1e",x"c0",x"87",x"f5"),
  1638 => (x"87",x"c6",x"fc",x"c0"),
  1639 => (x"ef",x"c0",x"49",x"70"),
  1640 => (x"ed",x"c3",x"87",x"e9"),
  1641 => (x"26",x"8e",x"f8",x"87"),
  1642 => (x"20",x"44",x"53",x"4f"),
  1643 => (x"6c",x"69",x"61",x"66"),
  1644 => (x"00",x"2e",x"64",x"65"),
  1645 => (x"74",x"6f",x"6f",x"42"),
  1646 => (x"2e",x"67",x"6e",x"69"),
  1647 => (x"1e",x"00",x"2e",x"2e"),
  1648 => (x"87",x"d4",x"e7",x"c0"),
  1649 => (x"87",x"f9",x"f2",x"c0"),
  1650 => (x"4f",x"26",x"87",x"f6"),
  1651 => (x"c8",x"f2",x"c2",x"1e"),
  1652 => (x"c2",x"78",x"c0",x"48"),
  1653 => (x"c0",x"48",x"f0",x"f1"),
  1654 => (x"87",x"fc",x"fd",x"78"),
  1655 => (x"48",x"c0",x"87",x"e1"),
  1656 => (x"00",x"00",x"4f",x"26"),
  1657 => (x"00",x"00",x"00",x"01"),
  1658 => (x"20",x"20",x"20",x"20"),
  1659 => (x"20",x"20",x"20",x"20"),
  1660 => (x"20",x"20",x"20",x"20"),
  1661 => (x"69",x"78",x"45",x"20"),
  1662 => (x"20",x"20",x"20",x"74"),
  1663 => (x"20",x"20",x"20",x"20"),
  1664 => (x"20",x"20",x"20",x"20"),
  1665 => (x"80",x"00",x"81",x"20"),
  1666 => (x"20",x"20",x"20",x"20"),
  1667 => (x"20",x"20",x"20",x"20"),
  1668 => (x"20",x"20",x"20",x"20"),
  1669 => (x"6b",x"63",x"61",x"42"),
  1670 => (x"00",x"12",x"d3",x"00"),
  1671 => (x"00",x"2c",x"9c",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"12",x"d3"),
  1674 => (x"00",x"00",x"2c",x"ba"),
  1675 => (x"d3",x"00",x"00",x"00"),
  1676 => (x"d8",x"00",x"00",x"12"),
  1677 => (x"00",x"00",x"00",x"2c"),
  1678 => (x"12",x"d3",x"00",x"00"),
  1679 => (x"2c",x"f6",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"12",x"d3",x"00"),
  1682 => (x"00",x"2d",x"14",x"00"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"00",x"00",x"12",x"d3"),
  1685 => (x"00",x"00",x"2d",x"32"),
  1686 => (x"d3",x"00",x"00",x"00"),
  1687 => (x"50",x"00",x"00",x"12"),
  1688 => (x"00",x"00",x"00",x"2d"),
  1689 => (x"12",x"d3",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"13",x"6e",x"00"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"00",x"00",x"00",x"00"),
  1695 => (x"48",x"f0",x"fe",x"1e"),
  1696 => (x"09",x"cd",x"78",x"c0"),
  1697 => (x"4f",x"26",x"09",x"79"),
  1698 => (x"f0",x"fe",x"1e",x"1e"),
  1699 => (x"26",x"48",x"7e",x"bf"),
  1700 => (x"fe",x"1e",x"4f",x"26"),
  1701 => (x"78",x"c1",x"48",x"f0"),
  1702 => (x"fe",x"1e",x"4f",x"26"),
  1703 => (x"78",x"c0",x"48",x"f0"),
  1704 => (x"71",x"1e",x"4f",x"26"),
  1705 => (x"52",x"52",x"c0",x"4a"),
  1706 => (x"5e",x"0e",x"4f",x"26"),
  1707 => (x"0e",x"5d",x"5c",x"5b"),
  1708 => (x"4d",x"71",x"86",x"f4"),
  1709 => (x"c1",x"7e",x"6d",x"97"),
  1710 => (x"6c",x"97",x"4c",x"a5"),
  1711 => (x"58",x"a6",x"c8",x"48"),
  1712 => (x"66",x"c4",x"48",x"6e"),
  1713 => (x"87",x"c5",x"05",x"a8"),
  1714 => (x"e6",x"c0",x"48",x"ff"),
  1715 => (x"87",x"ca",x"ff",x"87"),
  1716 => (x"97",x"49",x"a5",x"c2"),
  1717 => (x"a3",x"71",x"4b",x"6c"),
  1718 => (x"4b",x"6b",x"97",x"4b"),
  1719 => (x"6e",x"7e",x"6c",x"97"),
  1720 => (x"c8",x"80",x"c1",x"48"),
  1721 => (x"98",x"c7",x"58",x"a6"),
  1722 => (x"70",x"58",x"a6",x"cc"),
  1723 => (x"e1",x"fe",x"7c",x"97"),
  1724 => (x"f4",x"48",x"73",x"87"),
  1725 => (x"26",x"4d",x"26",x"8e"),
  1726 => (x"26",x"4b",x"26",x"4c"),
  1727 => (x"5b",x"5e",x"0e",x"4f"),
  1728 => (x"86",x"f4",x"0e",x"5c"),
  1729 => (x"66",x"d8",x"4c",x"71"),
  1730 => (x"9a",x"ff",x"c3",x"4a"),
  1731 => (x"97",x"4b",x"a4",x"c2"),
  1732 => (x"a1",x"73",x"49",x"6c"),
  1733 => (x"97",x"51",x"72",x"49"),
  1734 => (x"48",x"6e",x"7e",x"6c"),
  1735 => (x"a6",x"c8",x"80",x"c1"),
  1736 => (x"cc",x"98",x"c7",x"58"),
  1737 => (x"54",x"70",x"58",x"a6"),
  1738 => (x"ca",x"ff",x"8e",x"f4"),
  1739 => (x"fd",x"1e",x"1e",x"87"),
  1740 => (x"bf",x"e0",x"87",x"e8"),
  1741 => (x"e0",x"c0",x"49",x"4a"),
  1742 => (x"cb",x"02",x"99",x"c0"),
  1743 => (x"c2",x"1e",x"72",x"87"),
  1744 => (x"fe",x"49",x"ee",x"f5"),
  1745 => (x"86",x"c4",x"87",x"f7"),
  1746 => (x"70",x"87",x"fd",x"fc"),
  1747 => (x"87",x"c2",x"fd",x"7e"),
  1748 => (x"1e",x"4f",x"26",x"26"),
  1749 => (x"49",x"ee",x"f5",x"c2"),
  1750 => (x"c1",x"87",x"c7",x"fd"),
  1751 => (x"fc",x"49",x"ed",x"ec"),
  1752 => (x"f7",x"c3",x"87",x"da"),
  1753 => (x"0e",x"4f",x"26",x"87"),
  1754 => (x"5d",x"5c",x"5b",x"5e"),
  1755 => (x"c2",x"4d",x"71",x"0e"),
  1756 => (x"fc",x"49",x"ee",x"f5"),
  1757 => (x"4b",x"70",x"87",x"f4"),
  1758 => (x"04",x"ab",x"b7",x"c0"),
  1759 => (x"c3",x"87",x"c2",x"c3"),
  1760 => (x"c9",x"05",x"ab",x"f0"),
  1761 => (x"cb",x"f1",x"c1",x"87"),
  1762 => (x"c2",x"78",x"c1",x"48"),
  1763 => (x"e0",x"c3",x"87",x"e3"),
  1764 => (x"87",x"c9",x"05",x"ab"),
  1765 => (x"48",x"cf",x"f1",x"c1"),
  1766 => (x"d4",x"c2",x"78",x"c1"),
  1767 => (x"cf",x"f1",x"c1",x"87"),
  1768 => (x"87",x"c6",x"02",x"bf"),
  1769 => (x"4c",x"a3",x"c0",x"c2"),
  1770 => (x"4c",x"73",x"87",x"c2"),
  1771 => (x"bf",x"cb",x"f1",x"c1"),
  1772 => (x"87",x"e0",x"c0",x"02"),
  1773 => (x"b7",x"c4",x"49",x"74"),
  1774 => (x"f2",x"c1",x"91",x"29"),
  1775 => (x"4a",x"74",x"81",x"eb"),
  1776 => (x"92",x"c2",x"9a",x"cf"),
  1777 => (x"30",x"72",x"48",x"c1"),
  1778 => (x"ba",x"ff",x"4a",x"70"),
  1779 => (x"98",x"69",x"48",x"72"),
  1780 => (x"87",x"db",x"79",x"70"),
  1781 => (x"b7",x"c4",x"49",x"74"),
  1782 => (x"f2",x"c1",x"91",x"29"),
  1783 => (x"4a",x"74",x"81",x"eb"),
  1784 => (x"92",x"c2",x"9a",x"cf"),
  1785 => (x"30",x"72",x"48",x"c3"),
  1786 => (x"69",x"48",x"4a",x"70"),
  1787 => (x"75",x"79",x"70",x"b0"),
  1788 => (x"f0",x"c0",x"05",x"9d"),
  1789 => (x"48",x"d0",x"ff",x"87"),
  1790 => (x"ff",x"78",x"e1",x"c8"),
  1791 => (x"78",x"c5",x"48",x"d4"),
  1792 => (x"bf",x"cf",x"f1",x"c1"),
  1793 => (x"c3",x"87",x"c3",x"02"),
  1794 => (x"f1",x"c1",x"78",x"e0"),
  1795 => (x"c6",x"02",x"bf",x"cb"),
  1796 => (x"48",x"d4",x"ff",x"87"),
  1797 => (x"ff",x"78",x"f0",x"c3"),
  1798 => (x"78",x"73",x"48",x"d4"),
  1799 => (x"c8",x"48",x"d0",x"ff"),
  1800 => (x"e0",x"c0",x"78",x"e1"),
  1801 => (x"cf",x"f1",x"c1",x"78"),
  1802 => (x"c1",x"78",x"c0",x"48"),
  1803 => (x"c0",x"48",x"cb",x"f1"),
  1804 => (x"ee",x"f5",x"c2",x"78"),
  1805 => (x"87",x"f2",x"f9",x"49"),
  1806 => (x"b7",x"c0",x"4b",x"70"),
  1807 => (x"fe",x"fc",x"03",x"ab"),
  1808 => (x"26",x"48",x"c0",x"87"),
  1809 => (x"26",x"4c",x"26",x"4d"),
  1810 => (x"00",x"4f",x"26",x"4b"),
  1811 => (x"00",x"00",x"00",x"00"),
  1812 => (x"1e",x"00",x"00",x"00"),
  1813 => (x"fc",x"49",x"4a",x"71"),
  1814 => (x"4f",x"26",x"87",x"cd"),
  1815 => (x"72",x"4a",x"c0",x"1e"),
  1816 => (x"c1",x"91",x"c4",x"49"),
  1817 => (x"c0",x"81",x"eb",x"f2"),
  1818 => (x"d0",x"82",x"c1",x"79"),
  1819 => (x"ee",x"04",x"aa",x"b7"),
  1820 => (x"0e",x"4f",x"26",x"87"),
  1821 => (x"5d",x"5c",x"5b",x"5e"),
  1822 => (x"f8",x"4d",x"71",x"0e"),
  1823 => (x"4a",x"75",x"87",x"dc"),
  1824 => (x"92",x"2a",x"b7",x"c4"),
  1825 => (x"82",x"eb",x"f2",x"c1"),
  1826 => (x"9c",x"cf",x"4c",x"75"),
  1827 => (x"49",x"6a",x"94",x"c2"),
  1828 => (x"c3",x"2b",x"74",x"4b"),
  1829 => (x"74",x"48",x"c2",x"9b"),
  1830 => (x"ff",x"4c",x"70",x"30"),
  1831 => (x"71",x"48",x"74",x"bc"),
  1832 => (x"f7",x"7a",x"70",x"98"),
  1833 => (x"48",x"73",x"87",x"ec"),
  1834 => (x"00",x"87",x"d8",x"fe"),
  1835 => (x"70",x"00",x"00",x"00"),
  1836 => (x"70",x"70",x"70",x"70"),
  1837 => (x"70",x"70",x"70",x"70"),
  1838 => (x"70",x"70",x"70",x"70"),
  1839 => (x"70",x"70",x"70",x"70"),
  1840 => (x"70",x"70",x"70",x"70"),
  1841 => (x"70",x"70",x"70",x"70"),
  1842 => (x"70",x"70",x"70",x"70"),
  1843 => (x"70",x"70",x"70",x"70"),
  1844 => (x"70",x"70",x"70",x"70"),
  1845 => (x"70",x"70",x"70",x"70"),
  1846 => (x"70",x"70",x"70",x"70"),
  1847 => (x"70",x"70",x"70",x"70"),
  1848 => (x"70",x"70",x"70",x"70"),
  1849 => (x"70",x"70",x"70",x"70"),
  1850 => (x"1e",x"70",x"70",x"70"),
  1851 => (x"c8",x"48",x"d0",x"ff"),
  1852 => (x"48",x"71",x"78",x"e1"),
  1853 => (x"78",x"08",x"d4",x"ff"),
  1854 => (x"ff",x"1e",x"4f",x"26"),
  1855 => (x"e1",x"c8",x"48",x"d0"),
  1856 => (x"ff",x"48",x"71",x"78"),
  1857 => (x"c4",x"78",x"08",x"d4"),
  1858 => (x"d4",x"ff",x"48",x"66"),
  1859 => (x"4f",x"26",x"78",x"08"),
  1860 => (x"c4",x"4a",x"71",x"1e"),
  1861 => (x"72",x"1e",x"49",x"66"),
  1862 => (x"87",x"de",x"ff",x"49"),
  1863 => (x"c0",x"48",x"d0",x"ff"),
  1864 => (x"26",x"26",x"78",x"e0"),
  1865 => (x"1e",x"73",x"1e",x"4f"),
  1866 => (x"66",x"c8",x"4b",x"71"),
  1867 => (x"4a",x"73",x"1e",x"49"),
  1868 => (x"49",x"a2",x"e0",x"c1"),
  1869 => (x"26",x"87",x"d9",x"ff"),
  1870 => (x"4d",x"26",x"87",x"c4"),
  1871 => (x"4b",x"26",x"4c",x"26"),
  1872 => (x"73",x"1e",x"4f",x"26"),
  1873 => (x"4b",x"4a",x"71",x"1e"),
  1874 => (x"03",x"ab",x"b7",x"c2"),
  1875 => (x"49",x"a3",x"87",x"c8"),
  1876 => (x"9a",x"ff",x"c3",x"4a"),
  1877 => (x"a3",x"ce",x"87",x"c7"),
  1878 => (x"ff",x"c3",x"4a",x"49"),
  1879 => (x"49",x"66",x"c8",x"9a"),
  1880 => (x"fe",x"49",x"72",x"1e"),
  1881 => (x"ff",x"26",x"87",x"ea"),
  1882 => (x"ff",x"1e",x"87",x"d4"),
  1883 => (x"ff",x"c3",x"4a",x"d4"),
  1884 => (x"48",x"d0",x"ff",x"7a"),
  1885 => (x"de",x"78",x"e1",x"c0"),
  1886 => (x"f8",x"f5",x"c2",x"7a"),
  1887 => (x"48",x"49",x"7a",x"bf"),
  1888 => (x"7a",x"70",x"28",x"c8"),
  1889 => (x"28",x"d0",x"48",x"71"),
  1890 => (x"48",x"71",x"7a",x"70"),
  1891 => (x"7a",x"70",x"28",x"d8"),
  1892 => (x"c0",x"48",x"d0",x"ff"),
  1893 => (x"4f",x"26",x"78",x"e0"),
  1894 => (x"5c",x"5b",x"5e",x"0e"),
  1895 => (x"4c",x"71",x"0e",x"5d"),
  1896 => (x"bf",x"f8",x"f5",x"c2"),
  1897 => (x"29",x"74",x"49",x"4d"),
  1898 => (x"66",x"d0",x"4b",x"71"),
  1899 => (x"d4",x"83",x"c1",x"9b"),
  1900 => (x"04",x"ab",x"b7",x"66"),
  1901 => (x"4b",x"c0",x"87",x"c2"),
  1902 => (x"74",x"49",x"66",x"d0"),
  1903 => (x"75",x"b9",x"ff",x"31"),
  1904 => (x"74",x"4a",x"73",x"99"),
  1905 => (x"71",x"48",x"72",x"32"),
  1906 => (x"fc",x"f5",x"c2",x"b0"),
  1907 => (x"87",x"da",x"fe",x"58"),
  1908 => (x"4c",x"26",x"4d",x"26"),
  1909 => (x"4f",x"26",x"4b",x"26"),
  1910 => (x"48",x"d0",x"ff",x"1e"),
  1911 => (x"71",x"78",x"c9",x"c8"),
  1912 => (x"08",x"d4",x"ff",x"48"),
  1913 => (x"1e",x"4f",x"26",x"78"),
  1914 => (x"eb",x"49",x"4a",x"71"),
  1915 => (x"48",x"d0",x"ff",x"87"),
  1916 => (x"4f",x"26",x"78",x"c8"),
  1917 => (x"71",x"1e",x"73",x"1e"),
  1918 => (x"c8",x"f6",x"c2",x"4b"),
  1919 => (x"87",x"c3",x"02",x"bf"),
  1920 => (x"ff",x"87",x"eb",x"c2"),
  1921 => (x"c9",x"c8",x"48",x"d0"),
  1922 => (x"c0",x"49",x"73",x"78"),
  1923 => (x"d4",x"ff",x"b1",x"e0"),
  1924 => (x"c2",x"78",x"71",x"48"),
  1925 => (x"c0",x"48",x"fc",x"f5"),
  1926 => (x"02",x"66",x"c8",x"78"),
  1927 => (x"ff",x"c3",x"87",x"c5"),
  1928 => (x"c0",x"87",x"c2",x"49"),
  1929 => (x"c4",x"f6",x"c2",x"49"),
  1930 => (x"02",x"66",x"cc",x"59"),
  1931 => (x"d5",x"c5",x"87",x"c6"),
  1932 => (x"87",x"c4",x"4a",x"d5"),
  1933 => (x"4a",x"ff",x"ff",x"cf"),
  1934 => (x"5a",x"c8",x"f6",x"c2"),
  1935 => (x"48",x"c8",x"f6",x"c2"),
  1936 => (x"87",x"c4",x"78",x"c1"),
  1937 => (x"4c",x"26",x"4d",x"26"),
  1938 => (x"4f",x"26",x"4b",x"26"),
  1939 => (x"5c",x"5b",x"5e",x"0e"),
  1940 => (x"4a",x"71",x"0e",x"5d"),
  1941 => (x"bf",x"c4",x"f6",x"c2"),
  1942 => (x"02",x"9a",x"72",x"4c"),
  1943 => (x"c8",x"49",x"87",x"cb"),
  1944 => (x"ea",x"f7",x"c1",x"91"),
  1945 => (x"c4",x"83",x"71",x"4b"),
  1946 => (x"ea",x"fb",x"c1",x"87"),
  1947 => (x"13",x"4d",x"c0",x"4b"),
  1948 => (x"c2",x"99",x"74",x"49"),
  1949 => (x"b9",x"bf",x"c0",x"f6"),
  1950 => (x"71",x"48",x"d4",x"ff"),
  1951 => (x"2c",x"b7",x"c1",x"78"),
  1952 => (x"ad",x"b7",x"c8",x"85"),
  1953 => (x"c2",x"87",x"e8",x"04"),
  1954 => (x"48",x"bf",x"fc",x"f5"),
  1955 => (x"f6",x"c2",x"80",x"c8"),
  1956 => (x"ef",x"fe",x"58",x"c0"),
  1957 => (x"1e",x"73",x"1e",x"87"),
  1958 => (x"4a",x"13",x"4b",x"71"),
  1959 => (x"87",x"cb",x"02",x"9a"),
  1960 => (x"e7",x"fe",x"49",x"72"),
  1961 => (x"9a",x"4a",x"13",x"87"),
  1962 => (x"fe",x"87",x"f5",x"05"),
  1963 => (x"c2",x"1e",x"87",x"da"),
  1964 => (x"49",x"bf",x"fc",x"f5"),
  1965 => (x"48",x"fc",x"f5",x"c2"),
  1966 => (x"c4",x"78",x"a1",x"c1"),
  1967 => (x"03",x"a9",x"b7",x"c0"),
  1968 => (x"d4",x"ff",x"87",x"db"),
  1969 => (x"c0",x"f6",x"c2",x"48"),
  1970 => (x"f5",x"c2",x"78",x"bf"),
  1971 => (x"c2",x"49",x"bf",x"fc"),
  1972 => (x"c1",x"48",x"fc",x"f5"),
  1973 => (x"c0",x"c4",x"78",x"a1"),
  1974 => (x"e5",x"04",x"a9",x"b7"),
  1975 => (x"48",x"d0",x"ff",x"87"),
  1976 => (x"f6",x"c2",x"78",x"c8"),
  1977 => (x"78",x"c0",x"48",x"c8"),
  1978 => (x"00",x"00",x"4f",x"26"),
  1979 => (x"00",x"00",x"00",x"00"),
  1980 => (x"00",x"00",x"00",x"00"),
  1981 => (x"00",x"5f",x"5f",x"00"),
  1982 => (x"03",x"00",x"00",x"00"),
  1983 => (x"03",x"03",x"00",x"03"),
  1984 => (x"7f",x"14",x"00",x"00"),
  1985 => (x"7f",x"7f",x"14",x"7f"),
  1986 => (x"24",x"00",x"00",x"14"),
  1987 => (x"3a",x"6b",x"6b",x"2e"),
  1988 => (x"6a",x"4c",x"00",x"12"),
  1989 => (x"56",x"6c",x"18",x"36"),
  1990 => (x"7e",x"30",x"00",x"32"),
  1991 => (x"3a",x"77",x"59",x"4f"),
  1992 => (x"00",x"00",x"40",x"68"),
  1993 => (x"00",x"03",x"07",x"04"),
  1994 => (x"00",x"00",x"00",x"00"),
  1995 => (x"41",x"63",x"3e",x"1c"),
  1996 => (x"00",x"00",x"00",x"00"),
  1997 => (x"1c",x"3e",x"63",x"41"),
  1998 => (x"2a",x"08",x"00",x"00"),
  1999 => (x"3e",x"1c",x"1c",x"3e"),
  2000 => (x"08",x"00",x"08",x"2a"),
  2001 => (x"08",x"3e",x"3e",x"08"),
  2002 => (x"00",x"00",x"00",x"08"),
  2003 => (x"00",x"60",x"e0",x"80"),
  2004 => (x"08",x"00",x"00",x"00"),
  2005 => (x"08",x"08",x"08",x"08"),
  2006 => (x"00",x"00",x"00",x"08"),
  2007 => (x"00",x"60",x"60",x"00"),
  2008 => (x"60",x"40",x"00",x"00"),
  2009 => (x"06",x"0c",x"18",x"30"),
  2010 => (x"3e",x"00",x"01",x"03"),
  2011 => (x"7f",x"4d",x"59",x"7f"),
  2012 => (x"04",x"00",x"00",x"3e"),
  2013 => (x"00",x"7f",x"7f",x"06"),
  2014 => (x"42",x"00",x"00",x"00"),
  2015 => (x"4f",x"59",x"71",x"63"),
  2016 => (x"22",x"00",x"00",x"46"),
  2017 => (x"7f",x"49",x"49",x"63"),
  2018 => (x"1c",x"18",x"00",x"36"),
  2019 => (x"7f",x"7f",x"13",x"16"),
  2020 => (x"27",x"00",x"00",x"10"),
  2021 => (x"7d",x"45",x"45",x"67"),
  2022 => (x"3c",x"00",x"00",x"39"),
  2023 => (x"79",x"49",x"4b",x"7e"),
  2024 => (x"01",x"00",x"00",x"30"),
  2025 => (x"0f",x"79",x"71",x"01"),
  2026 => (x"36",x"00",x"00",x"07"),
  2027 => (x"7f",x"49",x"49",x"7f"),
  2028 => (x"06",x"00",x"00",x"36"),
  2029 => (x"3f",x"69",x"49",x"4f"),
  2030 => (x"00",x"00",x"00",x"1e"),
  2031 => (x"00",x"66",x"66",x"00"),
  2032 => (x"00",x"00",x"00",x"00"),
  2033 => (x"00",x"66",x"e6",x"80"),
  2034 => (x"08",x"00",x"00",x"00"),
  2035 => (x"22",x"14",x"14",x"08"),
  2036 => (x"14",x"00",x"00",x"22"),
  2037 => (x"14",x"14",x"14",x"14"),
  2038 => (x"22",x"00",x"00",x"14"),
  2039 => (x"08",x"14",x"14",x"22"),
  2040 => (x"02",x"00",x"00",x"08"),
  2041 => (x"0f",x"59",x"51",x"03"),
  2042 => (x"7f",x"3e",x"00",x"06"),
  2043 => (x"1f",x"55",x"5d",x"41"),
  2044 => (x"7e",x"00",x"00",x"1e"),
  2045 => (x"7f",x"09",x"09",x"7f"),
  2046 => (x"7f",x"00",x"00",x"7e"),
  2047 => (x"7f",x"49",x"49",x"7f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

