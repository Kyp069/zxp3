
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"40",x"7d",x"3d"),
     1 => (x"80",x"80",x"00",x"00"),
     2 => (x"00",x"7d",x"fd",x"80"),
     3 => (x"7f",x"7f",x"00",x"00"),
     4 => (x"44",x"6c",x"38",x"10"),
     5 => (x"00",x"00",x"00",x"00"),
     6 => (x"00",x"40",x"7f",x"3f"),
     7 => (x"0c",x"7c",x"7c",x"00"),
     8 => (x"78",x"7c",x"0c",x"18"),
     9 => (x"7c",x"7c",x"00",x"00"),
    10 => (x"78",x"7c",x"04",x"04"),
    11 => (x"7c",x"38",x"00",x"00"),
    12 => (x"38",x"7c",x"44",x"44"),
    13 => (x"fc",x"fc",x"00",x"00"),
    14 => (x"18",x"3c",x"24",x"24"),
    15 => (x"3c",x"18",x"00",x"00"),
    16 => (x"fc",x"fc",x"24",x"24"),
    17 => (x"7c",x"7c",x"00",x"00"),
    18 => (x"08",x"0c",x"04",x"04"),
    19 => (x"5c",x"48",x"00",x"00"),
    20 => (x"20",x"74",x"54",x"54"),
    21 => (x"3f",x"04",x"00",x"00"),
    22 => (x"00",x"44",x"44",x"7f"),
    23 => (x"7c",x"3c",x"00",x"00"),
    24 => (x"7c",x"7c",x"40",x"40"),
    25 => (x"3c",x"1c",x"00",x"00"),
    26 => (x"1c",x"3c",x"60",x"60"),
    27 => (x"60",x"7c",x"3c",x"00"),
    28 => (x"3c",x"7c",x"60",x"30"),
    29 => (x"38",x"6c",x"44",x"00"),
    30 => (x"44",x"6c",x"38",x"10"),
    31 => (x"bc",x"1c",x"00",x"00"),
    32 => (x"1c",x"3c",x"60",x"e0"),
    33 => (x"64",x"44",x"00",x"00"),
    34 => (x"44",x"4c",x"5c",x"74"),
    35 => (x"08",x"08",x"00",x"00"),
    36 => (x"41",x"41",x"77",x"3e"),
    37 => (x"00",x"00",x"00",x"00"),
    38 => (x"00",x"00",x"7f",x"7f"),
    39 => (x"41",x"41",x"00",x"00"),
    40 => (x"08",x"08",x"3e",x"77"),
    41 => (x"01",x"01",x"02",x"00"),
    42 => (x"01",x"02",x"02",x"03"),
    43 => (x"7f",x"7f",x"7f",x"00"),
    44 => (x"7f",x"7f",x"7f",x"7f"),
    45 => (x"1c",x"08",x"08",x"00"),
    46 => (x"7f",x"3e",x"3e",x"1c"),
    47 => (x"3e",x"7f",x"7f",x"7f"),
    48 => (x"08",x"1c",x"1c",x"3e"),
    49 => (x"18",x"10",x"00",x"08"),
    50 => (x"10",x"18",x"7c",x"7c"),
    51 => (x"30",x"10",x"00",x"00"),
    52 => (x"10",x"30",x"7c",x"7c"),
    53 => (x"60",x"30",x"10",x"00"),
    54 => (x"06",x"1e",x"78",x"60"),
    55 => (x"3c",x"66",x"42",x"00"),
    56 => (x"42",x"66",x"3c",x"18"),
    57 => (x"6a",x"38",x"78",x"00"),
    58 => (x"38",x"6c",x"c6",x"c2"),
    59 => (x"00",x"00",x"60",x"00"),
    60 => (x"60",x"00",x"00",x"60"),
    61 => (x"5b",x"5e",x"0e",x"00"),
    62 => (x"1e",x"0e",x"5d",x"5c"),
    63 => (x"ef",x"c2",x"4c",x"71"),
    64 => (x"c0",x"4d",x"bf",x"e9"),
    65 => (x"74",x"1e",x"c0",x"4b"),
    66 => (x"87",x"c7",x"02",x"ab"),
    67 => (x"c0",x"48",x"a6",x"c4"),
    68 => (x"c4",x"87",x"c5",x"78"),
    69 => (x"78",x"c1",x"48",x"a6"),
    70 => (x"73",x"1e",x"66",x"c4"),
    71 => (x"87",x"df",x"ee",x"49"),
    72 => (x"e0",x"c0",x"86",x"c8"),
    73 => (x"87",x"ef",x"ef",x"49"),
    74 => (x"6a",x"4a",x"a5",x"c4"),
    75 => (x"87",x"f0",x"f0",x"49"),
    76 => (x"cb",x"87",x"c6",x"f1"),
    77 => (x"c8",x"83",x"c1",x"85"),
    78 => (x"ff",x"04",x"ab",x"b7"),
    79 => (x"26",x"26",x"87",x"c7"),
    80 => (x"26",x"4c",x"26",x"4d"),
    81 => (x"1e",x"4f",x"26",x"4b"),
    82 => (x"ef",x"c2",x"4a",x"71"),
    83 => (x"ef",x"c2",x"5a",x"ed"),
    84 => (x"78",x"c7",x"48",x"ed"),
    85 => (x"87",x"dd",x"fe",x"49"),
    86 => (x"73",x"1e",x"4f",x"26"),
    87 => (x"c0",x"4a",x"71",x"1e"),
    88 => (x"d3",x"03",x"aa",x"b7"),
    89 => (x"eb",x"d2",x"c2",x"87"),
    90 => (x"87",x"c4",x"05",x"bf"),
    91 => (x"87",x"c2",x"4b",x"c1"),
    92 => (x"d2",x"c2",x"4b",x"c0"),
    93 => (x"87",x"c4",x"5b",x"ef"),
    94 => (x"5a",x"ef",x"d2",x"c2"),
    95 => (x"bf",x"eb",x"d2",x"c2"),
    96 => (x"c1",x"9a",x"c1",x"4a"),
    97 => (x"ec",x"49",x"a2",x"c0"),
    98 => (x"48",x"fc",x"87",x"e8"),
    99 => (x"bf",x"eb",x"d2",x"c2"),
   100 => (x"87",x"ef",x"fe",x"78"),
   101 => (x"c4",x"4a",x"71",x"1e"),
   102 => (x"49",x"72",x"1e",x"66"),
   103 => (x"26",x"87",x"ee",x"e9"),
   104 => (x"c2",x"1e",x"4f",x"26"),
   105 => (x"49",x"bf",x"eb",x"d2"),
   106 => (x"c2",x"87",x"f3",x"e5"),
   107 => (x"e8",x"48",x"e1",x"ef"),
   108 => (x"ef",x"c2",x"78",x"bf"),
   109 => (x"bf",x"ec",x"48",x"dd"),
   110 => (x"e1",x"ef",x"c2",x"78"),
   111 => (x"c3",x"49",x"4a",x"bf"),
   112 => (x"b7",x"c8",x"99",x"ff"),
   113 => (x"71",x"48",x"72",x"2a"),
   114 => (x"e9",x"ef",x"c2",x"b0"),
   115 => (x"0e",x"4f",x"26",x"58"),
   116 => (x"5d",x"5c",x"5b",x"5e"),
   117 => (x"ff",x"4b",x"71",x"0e"),
   118 => (x"ef",x"c2",x"87",x"c8"),
   119 => (x"50",x"c0",x"48",x"dc"),
   120 => (x"d9",x"e5",x"49",x"73"),
   121 => (x"4c",x"49",x"70",x"87"),
   122 => (x"ee",x"cb",x"9c",x"c2"),
   123 => (x"87",x"c3",x"cb",x"49"),
   124 => (x"c2",x"4d",x"49",x"70"),
   125 => (x"bf",x"97",x"dc",x"ef"),
   126 => (x"87",x"e2",x"c1",x"05"),
   127 => (x"c2",x"49",x"66",x"d0"),
   128 => (x"99",x"bf",x"e5",x"ef"),
   129 => (x"d4",x"87",x"d6",x"05"),
   130 => (x"ef",x"c2",x"49",x"66"),
   131 => (x"05",x"99",x"bf",x"dd"),
   132 => (x"49",x"73",x"87",x"cb"),
   133 => (x"70",x"87",x"e7",x"e4"),
   134 => (x"c1",x"c1",x"02",x"98"),
   135 => (x"fe",x"4c",x"c1",x"87"),
   136 => (x"49",x"75",x"87",x"c0"),
   137 => (x"70",x"87",x"d8",x"ca"),
   138 => (x"87",x"c6",x"02",x"98"),
   139 => (x"48",x"dc",x"ef",x"c2"),
   140 => (x"ef",x"c2",x"50",x"c1"),
   141 => (x"05",x"bf",x"97",x"dc"),
   142 => (x"c2",x"87",x"e3",x"c0"),
   143 => (x"49",x"bf",x"e5",x"ef"),
   144 => (x"05",x"99",x"66",x"d0"),
   145 => (x"c2",x"87",x"d6",x"ff"),
   146 => (x"49",x"bf",x"dd",x"ef"),
   147 => (x"05",x"99",x"66",x"d4"),
   148 => (x"73",x"87",x"ca",x"ff"),
   149 => (x"87",x"e6",x"e3",x"49"),
   150 => (x"fe",x"05",x"98",x"70"),
   151 => (x"48",x"74",x"87",x"ff"),
   152 => (x"0e",x"87",x"dc",x"fb"),
   153 => (x"5d",x"5c",x"5b",x"5e"),
   154 => (x"c0",x"86",x"f4",x"0e"),
   155 => (x"bf",x"ec",x"4c",x"4d"),
   156 => (x"48",x"a6",x"c4",x"7e"),
   157 => (x"bf",x"e9",x"ef",x"c2"),
   158 => (x"c0",x"1e",x"c1",x"78"),
   159 => (x"fd",x"49",x"c7",x"1e"),
   160 => (x"86",x"c8",x"87",x"cd"),
   161 => (x"cd",x"02",x"98",x"70"),
   162 => (x"fb",x"49",x"ff",x"87"),
   163 => (x"da",x"c1",x"87",x"cc"),
   164 => (x"87",x"ea",x"e2",x"49"),
   165 => (x"ef",x"c2",x"4d",x"c1"),
   166 => (x"02",x"bf",x"97",x"dc"),
   167 => (x"fc",x"cf",x"87",x"c3"),
   168 => (x"e1",x"ef",x"c2",x"87"),
   169 => (x"d2",x"c2",x"4b",x"bf"),
   170 => (x"c0",x"05",x"bf",x"eb"),
   171 => (x"fd",x"c3",x"87",x"e9"),
   172 => (x"87",x"ca",x"e2",x"49"),
   173 => (x"e2",x"49",x"fa",x"c3"),
   174 => (x"49",x"73",x"87",x"c4"),
   175 => (x"71",x"99",x"ff",x"c3"),
   176 => (x"fb",x"49",x"c0",x"1e"),
   177 => (x"49",x"73",x"87",x"ce"),
   178 => (x"71",x"29",x"b7",x"c8"),
   179 => (x"fb",x"49",x"c1",x"1e"),
   180 => (x"86",x"c8",x"87",x"c2"),
   181 => (x"c2",x"87",x"fa",x"c5"),
   182 => (x"4b",x"bf",x"e5",x"ef"),
   183 => (x"87",x"dd",x"02",x"9b"),
   184 => (x"bf",x"e7",x"d2",x"c2"),
   185 => (x"87",x"d7",x"c7",x"49"),
   186 => (x"c4",x"05",x"98",x"70"),
   187 => (x"d2",x"4b",x"c0",x"87"),
   188 => (x"49",x"e0",x"c2",x"87"),
   189 => (x"c2",x"87",x"fc",x"c6"),
   190 => (x"c6",x"58",x"eb",x"d2"),
   191 => (x"e7",x"d2",x"c2",x"87"),
   192 => (x"73",x"78",x"c0",x"48"),
   193 => (x"05",x"99",x"c2",x"49"),
   194 => (x"eb",x"c3",x"87",x"cd"),
   195 => (x"87",x"ee",x"e0",x"49"),
   196 => (x"99",x"c2",x"49",x"70"),
   197 => (x"fb",x"87",x"c2",x"02"),
   198 => (x"c1",x"49",x"73",x"4c"),
   199 => (x"87",x"cd",x"05",x"99"),
   200 => (x"e0",x"49",x"f4",x"c3"),
   201 => (x"49",x"70",x"87",x"d8"),
   202 => (x"c2",x"02",x"99",x"c2"),
   203 => (x"73",x"4c",x"fa",x"87"),
   204 => (x"05",x"99",x"c8",x"49"),
   205 => (x"f5",x"c3",x"87",x"cd"),
   206 => (x"87",x"c2",x"e0",x"49"),
   207 => (x"99",x"c2",x"49",x"70"),
   208 => (x"c2",x"87",x"d4",x"02"),
   209 => (x"02",x"bf",x"ed",x"ef"),
   210 => (x"c1",x"48",x"87",x"c9"),
   211 => (x"f1",x"ef",x"c2",x"88"),
   212 => (x"ff",x"87",x"c2",x"58"),
   213 => (x"73",x"4d",x"c1",x"4c"),
   214 => (x"05",x"99",x"c4",x"49"),
   215 => (x"f2",x"c3",x"87",x"ce"),
   216 => (x"d9",x"df",x"ff",x"49"),
   217 => (x"c2",x"49",x"70",x"87"),
   218 => (x"87",x"db",x"02",x"99"),
   219 => (x"bf",x"ed",x"ef",x"c2"),
   220 => (x"b7",x"c7",x"48",x"7e"),
   221 => (x"87",x"cb",x"03",x"a8"),
   222 => (x"80",x"c1",x"48",x"6e"),
   223 => (x"58",x"f1",x"ef",x"c2"),
   224 => (x"fe",x"87",x"c2",x"c0"),
   225 => (x"c3",x"4d",x"c1",x"4c"),
   226 => (x"de",x"ff",x"49",x"fd"),
   227 => (x"49",x"70",x"87",x"f0"),
   228 => (x"d5",x"02",x"99",x"c2"),
   229 => (x"ed",x"ef",x"c2",x"87"),
   230 => (x"c9",x"c0",x"02",x"bf"),
   231 => (x"ed",x"ef",x"c2",x"87"),
   232 => (x"c0",x"78",x"c0",x"48"),
   233 => (x"4c",x"fd",x"87",x"c2"),
   234 => (x"fa",x"c3",x"4d",x"c1"),
   235 => (x"cd",x"de",x"ff",x"49"),
   236 => (x"c2",x"49",x"70",x"87"),
   237 => (x"87",x"d9",x"02",x"99"),
   238 => (x"bf",x"ed",x"ef",x"c2"),
   239 => (x"a8",x"b7",x"c7",x"48"),
   240 => (x"87",x"c9",x"c0",x"03"),
   241 => (x"48",x"ed",x"ef",x"c2"),
   242 => (x"c2",x"c0",x"78",x"c7"),
   243 => (x"c1",x"4c",x"fc",x"87"),
   244 => (x"ac",x"b7",x"c0",x"4d"),
   245 => (x"87",x"d1",x"c0",x"03"),
   246 => (x"c1",x"4a",x"66",x"c4"),
   247 => (x"02",x"6a",x"82",x"d8"),
   248 => (x"6a",x"87",x"c6",x"c0"),
   249 => (x"73",x"49",x"74",x"4b"),
   250 => (x"c3",x"1e",x"c0",x"0f"),
   251 => (x"da",x"c1",x"1e",x"f0"),
   252 => (x"87",x"db",x"f7",x"49"),
   253 => (x"98",x"70",x"86",x"c8"),
   254 => (x"87",x"e2",x"c0",x"02"),
   255 => (x"c2",x"48",x"a6",x"c8"),
   256 => (x"78",x"bf",x"ed",x"ef"),
   257 => (x"cb",x"49",x"66",x"c8"),
   258 => (x"48",x"66",x"c4",x"91"),
   259 => (x"7e",x"70",x"80",x"71"),
   260 => (x"c0",x"02",x"bf",x"6e"),
   261 => (x"bf",x"6e",x"87",x"c8"),
   262 => (x"49",x"66",x"c8",x"4b"),
   263 => (x"9d",x"75",x"0f",x"73"),
   264 => (x"87",x"c8",x"c0",x"02"),
   265 => (x"bf",x"ed",x"ef",x"c2"),
   266 => (x"87",x"c9",x"f3",x"49"),
   267 => (x"bf",x"ef",x"d2",x"c2"),
   268 => (x"87",x"dd",x"c0",x"02"),
   269 => (x"87",x"c7",x"c2",x"49"),
   270 => (x"c0",x"02",x"98",x"70"),
   271 => (x"ef",x"c2",x"87",x"d3"),
   272 => (x"f2",x"49",x"bf",x"ed"),
   273 => (x"49",x"c0",x"87",x"ef"),
   274 => (x"c2",x"87",x"cf",x"f4"),
   275 => (x"c0",x"48",x"ef",x"d2"),
   276 => (x"f3",x"8e",x"f4",x"78"),
   277 => (x"5e",x"0e",x"87",x"e9"),
   278 => (x"0e",x"5d",x"5c",x"5b"),
   279 => (x"c2",x"4c",x"71",x"1e"),
   280 => (x"49",x"bf",x"e9",x"ef"),
   281 => (x"4d",x"a1",x"cd",x"c1"),
   282 => (x"69",x"81",x"d1",x"c1"),
   283 => (x"02",x"9c",x"74",x"7e"),
   284 => (x"a5",x"c4",x"87",x"cf"),
   285 => (x"c2",x"7b",x"74",x"4b"),
   286 => (x"49",x"bf",x"e9",x"ef"),
   287 => (x"6e",x"87",x"c8",x"f3"),
   288 => (x"05",x"9c",x"74",x"7b"),
   289 => (x"4b",x"c0",x"87",x"c4"),
   290 => (x"4b",x"c1",x"87",x"c2"),
   291 => (x"c9",x"f3",x"49",x"73"),
   292 => (x"02",x"66",x"d4",x"87"),
   293 => (x"da",x"49",x"87",x"c7"),
   294 => (x"c2",x"4a",x"70",x"87"),
   295 => (x"c2",x"4a",x"c0",x"87"),
   296 => (x"26",x"5a",x"f3",x"d2"),
   297 => (x"00",x"87",x"d8",x"f2"),
   298 => (x"00",x"00",x"00",x"00"),
   299 => (x"00",x"00",x"00",x"00"),
   300 => (x"1e",x"00",x"00",x"00"),
   301 => (x"c8",x"ff",x"4a",x"71"),
   302 => (x"a1",x"72",x"49",x"bf"),
   303 => (x"1e",x"4f",x"26",x"48"),
   304 => (x"89",x"bf",x"c8",x"ff"),
   305 => (x"c0",x"c0",x"c0",x"c2"),
   306 => (x"01",x"a9",x"c0",x"c0"),
   307 => (x"4a",x"c0",x"87",x"c4"),
   308 => (x"4a",x"c1",x"87",x"c2"),
   309 => (x"4f",x"26",x"48",x"72"),
   310 => (x"5c",x"5b",x"5e",x"0e"),
   311 => (x"4b",x"71",x"0e",x"5d"),
   312 => (x"d0",x"4c",x"d4",x"ff"),
   313 => (x"78",x"c0",x"48",x"66"),
   314 => (x"db",x"ff",x"49",x"d6"),
   315 => (x"ff",x"c3",x"87",x"c8"),
   316 => (x"c3",x"49",x"6c",x"7c"),
   317 => (x"4d",x"71",x"99",x"ff"),
   318 => (x"99",x"f0",x"c3",x"49"),
   319 => (x"05",x"a9",x"e0",x"c1"),
   320 => (x"ff",x"c3",x"87",x"cb"),
   321 => (x"c3",x"48",x"6c",x"7c"),
   322 => (x"08",x"66",x"d0",x"98"),
   323 => (x"7c",x"ff",x"c3",x"78"),
   324 => (x"c8",x"49",x"4a",x"6c"),
   325 => (x"7c",x"ff",x"c3",x"31"),
   326 => (x"b2",x"71",x"4a",x"6c"),
   327 => (x"31",x"c8",x"49",x"72"),
   328 => (x"6c",x"7c",x"ff",x"c3"),
   329 => (x"72",x"b2",x"71",x"4a"),
   330 => (x"c3",x"31",x"c8",x"49"),
   331 => (x"4a",x"6c",x"7c",x"ff"),
   332 => (x"d0",x"ff",x"b2",x"71"),
   333 => (x"78",x"e0",x"c0",x"48"),
   334 => (x"c2",x"02",x"9b",x"73"),
   335 => (x"75",x"7b",x"72",x"87"),
   336 => (x"26",x"4d",x"26",x"48"),
   337 => (x"26",x"4b",x"26",x"4c"),
   338 => (x"4f",x"26",x"1e",x"4f"),
   339 => (x"5c",x"5b",x"5e",x"0e"),
   340 => (x"76",x"86",x"f8",x"0e"),
   341 => (x"49",x"a6",x"c8",x"1e"),
   342 => (x"c4",x"87",x"fd",x"fd"),
   343 => (x"6e",x"4b",x"70",x"86"),
   344 => (x"03",x"a8",x"c3",x"48"),
   345 => (x"73",x"87",x"f0",x"c2"),
   346 => (x"9a",x"f0",x"c3",x"4a"),
   347 => (x"02",x"aa",x"d0",x"c1"),
   348 => (x"e0",x"c1",x"87",x"c7"),
   349 => (x"de",x"c2",x"05",x"aa"),
   350 => (x"c8",x"49",x"73",x"87"),
   351 => (x"87",x"c3",x"02",x"99"),
   352 => (x"73",x"87",x"c6",x"ff"),
   353 => (x"c2",x"9c",x"c3",x"4c"),
   354 => (x"c2",x"c1",x"05",x"ac"),
   355 => (x"49",x"66",x"c4",x"87"),
   356 => (x"1e",x"71",x"31",x"c9"),
   357 => (x"d4",x"4a",x"66",x"c4"),
   358 => (x"f1",x"ef",x"c2",x"92"),
   359 => (x"fe",x"81",x"72",x"49"),
   360 => (x"d8",x"87",x"ef",x"d0"),
   361 => (x"cd",x"d8",x"ff",x"49"),
   362 => (x"1e",x"c0",x"c8",x"87"),
   363 => (x"49",x"ce",x"de",x"c2"),
   364 => (x"87",x"eb",x"ec",x"fd"),
   365 => (x"c0",x"48",x"d0",x"ff"),
   366 => (x"de",x"c2",x"78",x"e0"),
   367 => (x"66",x"cc",x"1e",x"ce"),
   368 => (x"c2",x"92",x"d4",x"4a"),
   369 => (x"72",x"49",x"f1",x"ef"),
   370 => (x"f6",x"ce",x"fe",x"81"),
   371 => (x"c1",x"86",x"cc",x"87"),
   372 => (x"c2",x"c1",x"05",x"ac"),
   373 => (x"49",x"66",x"c4",x"87"),
   374 => (x"1e",x"71",x"31",x"c9"),
   375 => (x"d4",x"4a",x"66",x"c4"),
   376 => (x"f1",x"ef",x"c2",x"92"),
   377 => (x"fe",x"81",x"72",x"49"),
   378 => (x"c2",x"87",x"e7",x"cf"),
   379 => (x"c8",x"1e",x"ce",x"de"),
   380 => (x"92",x"d4",x"4a",x"66"),
   381 => (x"49",x"f1",x"ef",x"c2"),
   382 => (x"cc",x"fe",x"81",x"72"),
   383 => (x"49",x"d7",x"87",x"f6"),
   384 => (x"87",x"f2",x"d6",x"ff"),
   385 => (x"c2",x"1e",x"c0",x"c8"),
   386 => (x"fd",x"49",x"ce",x"de"),
   387 => (x"cc",x"87",x"e9",x"ea"),
   388 => (x"48",x"d0",x"ff",x"86"),
   389 => (x"f8",x"78",x"e0",x"c0"),
   390 => (x"87",x"e7",x"fc",x"8e"),
   391 => (x"5c",x"5b",x"5e",x"0e"),
   392 => (x"71",x"1e",x"0e",x"5d"),
   393 => (x"4c",x"d4",x"ff",x"4d"),
   394 => (x"48",x"7e",x"66",x"d4"),
   395 => (x"06",x"a8",x"b7",x"c3"),
   396 => (x"48",x"c0",x"87",x"c5"),
   397 => (x"75",x"87",x"e2",x"c1"),
   398 => (x"e2",x"dd",x"fe",x"49"),
   399 => (x"c4",x"1e",x"75",x"87"),
   400 => (x"93",x"d4",x"4b",x"66"),
   401 => (x"83",x"f1",x"ef",x"c2"),
   402 => (x"c6",x"fe",x"49",x"73"),
   403 => (x"83",x"c8",x"87",x"f3"),
   404 => (x"d0",x"ff",x"4b",x"6b"),
   405 => (x"78",x"e1",x"c8",x"48"),
   406 => (x"49",x"73",x"7c",x"dd"),
   407 => (x"71",x"99",x"ff",x"c3"),
   408 => (x"c8",x"49",x"73",x"7c"),
   409 => (x"ff",x"c3",x"29",x"b7"),
   410 => (x"73",x"7c",x"71",x"99"),
   411 => (x"29",x"b7",x"d0",x"49"),
   412 => (x"71",x"99",x"ff",x"c3"),
   413 => (x"d8",x"49",x"73",x"7c"),
   414 => (x"7c",x"71",x"29",x"b7"),
   415 => (x"7c",x"7c",x"7c",x"c0"),
   416 => (x"7c",x"7c",x"7c",x"7c"),
   417 => (x"7c",x"7c",x"7c",x"7c"),
   418 => (x"78",x"e0",x"c0",x"7c"),
   419 => (x"dc",x"1e",x"66",x"c4"),
   420 => (x"c6",x"d5",x"ff",x"49"),
   421 => (x"73",x"86",x"c8",x"87"),
   422 => (x"e4",x"fa",x"26",x"48"),
   423 => (x"db",x"c2",x"1e",x"87"),
   424 => (x"c1",x"49",x"bf",x"c6"),
   425 => (x"ca",x"db",x"c2",x"b9"),
   426 => (x"48",x"d4",x"ff",x"59"),
   427 => (x"ff",x"78",x"ff",x"c3"),
   428 => (x"e1",x"c0",x"48",x"d0"),
   429 => (x"48",x"d4",x"ff",x"78"),
   430 => (x"31",x"c4",x"78",x"c1"),
   431 => (x"d0",x"ff",x"78",x"71"),
   432 => (x"78",x"e0",x"c0",x"48"),
   433 => (x"00",x"00",x"4f",x"26"),
   434 => (x"c1",x"1e",x"00",x"00"),
   435 => (x"c0",x"48",x"d0",x"e3"),
   436 => (x"d6",x"dc",x"c2",x"50"),
   437 => (x"de",x"fe",x"49",x"bf"),
   438 => (x"e3",x"c1",x"87",x"eb"),
   439 => (x"50",x"c1",x"48",x"d0"),
   440 => (x"bf",x"da",x"dc",x"c2"),
   441 => (x"dc",x"de",x"fe",x"49"),
   442 => (x"d0",x"e3",x"c1",x"87"),
   443 => (x"c2",x"50",x"c2",x"48"),
   444 => (x"49",x"bf",x"de",x"dc"),
   445 => (x"87",x"cd",x"de",x"fe"),
   446 => (x"48",x"d0",x"e3",x"c1"),
   447 => (x"dc",x"c2",x"50",x"c3"),
   448 => (x"fe",x"49",x"bf",x"e2"),
   449 => (x"c0",x"87",x"fe",x"dd"),
   450 => (x"e6",x"dc",x"c2",x"1e"),
   451 => (x"cb",x"fc",x"49",x"bf"),
   452 => (x"26",x"48",x"c0",x"87"),
   453 => (x"27",x"2a",x"4f",x"26"),
   454 => (x"27",x"36",x"00",x"00"),
   455 => (x"27",x"42",x"00",x"00"),
   456 => (x"27",x"4e",x"00",x"00"),
   457 => (x"27",x"5a",x"00",x"00"),
   458 => (x"30",x"30",x"00",x"00"),
   459 => (x"20",x"20",x"20",x"20"),
   460 => (x"43",x"53",x"20",x"20"),
   461 => (x"31",x"30",x"00",x"52"),
   462 => (x"20",x"20",x"20",x"20"),
   463 => (x"43",x"53",x"20",x"20"),
   464 => (x"32",x"30",x"00",x"52"),
   465 => (x"20",x"20",x"20",x"20"),
   466 => (x"43",x"53",x"20",x"20"),
   467 => (x"33",x"30",x"00",x"52"),
   468 => (x"20",x"20",x"20",x"20"),
   469 => (x"43",x"53",x"20",x"20"),
   470 => (x"58",x"5a",x"00",x"52"),
   471 => (x"20",x"20",x"33",x"50"),
   472 => (x"48",x"56",x"20",x"20"),
   473 => (x"48",x"56",x"00",x"44"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

