
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"f0",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"f0",x"f0",x"c2"),
    14 => (x"48",x"e8",x"dd",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ef",x"e1"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d4",x"02",x"99",x"71"),
    50 => (x"ff",x"48",x"12",x"87"),
    51 => (x"c4",x"78",x"08",x"d4"),
    52 => (x"c1",x"48",x"49",x"66"),
    53 => (x"58",x"a6",x"c8",x"88"),
    54 => (x"ec",x"05",x"99",x"71"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"66",x"c4",x"4a",x"71"),
    57 => (x"88",x"c1",x"48",x"49"),
    58 => (x"71",x"58",x"a6",x"c8"),
    59 => (x"87",x"d6",x"02",x"99"),
    60 => (x"c3",x"48",x"d4",x"ff"),
    61 => (x"52",x"68",x"78",x"ff"),
    62 => (x"48",x"49",x"66",x"c4"),
    63 => (x"a6",x"c8",x"88",x"c1"),
    64 => (x"05",x"99",x"71",x"58"),
    65 => (x"4f",x"26",x"87",x"ea"),
    66 => (x"ff",x"1e",x"73",x"1e"),
    67 => (x"ff",x"c3",x"4b",x"d4"),
    68 => (x"c3",x"4a",x"6b",x"7b"),
    69 => (x"49",x"6b",x"7b",x"ff"),
    70 => (x"b1",x"72",x"32",x"c8"),
    71 => (x"6b",x"7b",x"ff",x"c3"),
    72 => (x"71",x"31",x"c8",x"4a"),
    73 => (x"7b",x"ff",x"c3",x"b2"),
    74 => (x"32",x"c8",x"49",x"6b"),
    75 => (x"48",x"71",x"b1",x"72"),
    76 => (x"4d",x"26",x"87",x"c4"),
    77 => (x"4b",x"26",x"4c",x"26"),
    78 => (x"5e",x"0e",x"4f",x"26"),
    79 => (x"0e",x"5d",x"5c",x"5b"),
    80 => (x"d4",x"ff",x"4a",x"71"),
    81 => (x"c3",x"49",x"72",x"4c"),
    82 => (x"7c",x"71",x"99",x"ff"),
    83 => (x"bf",x"e8",x"dd",x"c2"),
    84 => (x"d0",x"87",x"c8",x"05"),
    85 => (x"30",x"c9",x"48",x"66"),
    86 => (x"d0",x"58",x"a6",x"d4"),
    87 => (x"29",x"d8",x"49",x"66"),
    88 => (x"71",x"99",x"ff",x"c3"),
    89 => (x"49",x"66",x"d0",x"7c"),
    90 => (x"ff",x"c3",x"29",x"d0"),
    91 => (x"d0",x"7c",x"71",x"99"),
    92 => (x"29",x"c8",x"49",x"66"),
    93 => (x"71",x"99",x"ff",x"c3"),
    94 => (x"49",x"66",x"d0",x"7c"),
    95 => (x"71",x"99",x"ff",x"c3"),
    96 => (x"d0",x"49",x"72",x"7c"),
    97 => (x"99",x"ff",x"c3",x"29"),
    98 => (x"4b",x"6c",x"7c",x"71"),
    99 => (x"4d",x"ff",x"f0",x"c9"),
   100 => (x"05",x"ab",x"ff",x"c3"),
   101 => (x"ff",x"c3",x"87",x"d0"),
   102 => (x"c1",x"4b",x"6c",x"7c"),
   103 => (x"87",x"c6",x"02",x"8d"),
   104 => (x"02",x"ab",x"ff",x"c3"),
   105 => (x"48",x"73",x"87",x"f0"),
   106 => (x"1e",x"87",x"c7",x"fe"),
   107 => (x"d4",x"ff",x"49",x"c0"),
   108 => (x"78",x"ff",x"c3",x"48"),
   109 => (x"c8",x"c3",x"81",x"c1"),
   110 => (x"f1",x"04",x"a9",x"b7"),
   111 => (x"1e",x"4f",x"26",x"87"),
   112 => (x"87",x"e7",x"1e",x"73"),
   113 => (x"4b",x"df",x"f8",x"c4"),
   114 => (x"ff",x"c0",x"1e",x"c0"),
   115 => (x"49",x"f7",x"c1",x"f0"),
   116 => (x"c4",x"87",x"e7",x"fd"),
   117 => (x"05",x"a8",x"c1",x"86"),
   118 => (x"ff",x"87",x"ea",x"c0"),
   119 => (x"ff",x"c3",x"48",x"d4"),
   120 => (x"c0",x"c0",x"c1",x"78"),
   121 => (x"1e",x"c0",x"c0",x"c0"),
   122 => (x"c1",x"f0",x"e1",x"c0"),
   123 => (x"c9",x"fd",x"49",x"e9"),
   124 => (x"70",x"86",x"c4",x"87"),
   125 => (x"87",x"ca",x"05",x"98"),
   126 => (x"c3",x"48",x"d4",x"ff"),
   127 => (x"48",x"c1",x"78",x"ff"),
   128 => (x"e6",x"fe",x"87",x"cb"),
   129 => (x"05",x"8b",x"c1",x"87"),
   130 => (x"c0",x"87",x"fd",x"fe"),
   131 => (x"87",x"e6",x"fc",x"48"),
   132 => (x"ff",x"1e",x"73",x"1e"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"c0",x"4b",x"d3",x"78"),
   135 => (x"f0",x"ff",x"c0",x"1e"),
   136 => (x"fc",x"49",x"c1",x"c1"),
   137 => (x"86",x"c4",x"87",x"d4"),
   138 => (x"ca",x"05",x"98",x"70"),
   139 => (x"48",x"d4",x"ff",x"87"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"fd",x"87",x"cb",x"48"),
   142 => (x"8b",x"c1",x"87",x"f1"),
   143 => (x"87",x"db",x"ff",x"05"),
   144 => (x"f1",x"fb",x"48",x"c0"),
   145 => (x"5b",x"5e",x"0e",x"87"),
   146 => (x"d4",x"ff",x"0e",x"5c"),
   147 => (x"87",x"db",x"fd",x"4c"),
   148 => (x"c0",x"1e",x"ea",x"c6"),
   149 => (x"c8",x"c1",x"f0",x"e1"),
   150 => (x"87",x"de",x"fb",x"49"),
   151 => (x"a8",x"c1",x"86",x"c4"),
   152 => (x"fe",x"87",x"c8",x"02"),
   153 => (x"48",x"c0",x"87",x"ea"),
   154 => (x"fa",x"87",x"e2",x"c1"),
   155 => (x"49",x"70",x"87",x"da"),
   156 => (x"99",x"ff",x"ff",x"cf"),
   157 => (x"02",x"a9",x"ea",x"c6"),
   158 => (x"d3",x"fe",x"87",x"c8"),
   159 => (x"c1",x"48",x"c0",x"87"),
   160 => (x"ff",x"c3",x"87",x"cb"),
   161 => (x"4b",x"f1",x"c0",x"7c"),
   162 => (x"70",x"87",x"f4",x"fc"),
   163 => (x"eb",x"c0",x"02",x"98"),
   164 => (x"c0",x"1e",x"c0",x"87"),
   165 => (x"fa",x"c1",x"f0",x"ff"),
   166 => (x"87",x"de",x"fa",x"49"),
   167 => (x"98",x"70",x"86",x"c4"),
   168 => (x"c3",x"87",x"d9",x"05"),
   169 => (x"49",x"6c",x"7c",x"ff"),
   170 => (x"7c",x"7c",x"ff",x"c3"),
   171 => (x"c0",x"c1",x"7c",x"7c"),
   172 => (x"87",x"c4",x"02",x"99"),
   173 => (x"87",x"d5",x"48",x"c1"),
   174 => (x"87",x"d1",x"48",x"c0"),
   175 => (x"c4",x"05",x"ab",x"c2"),
   176 => (x"c8",x"48",x"c0",x"87"),
   177 => (x"05",x"8b",x"c1",x"87"),
   178 => (x"c0",x"87",x"fd",x"fe"),
   179 => (x"87",x"e4",x"f9",x"48"),
   180 => (x"c2",x"1e",x"73",x"1e"),
   181 => (x"c1",x"48",x"e8",x"dd"),
   182 => (x"ff",x"4b",x"c7",x"78"),
   183 => (x"78",x"c2",x"48",x"d0"),
   184 => (x"ff",x"87",x"c8",x"fb"),
   185 => (x"78",x"c3",x"48",x"d0"),
   186 => (x"e5",x"c0",x"1e",x"c0"),
   187 => (x"49",x"c0",x"c1",x"d0"),
   188 => (x"c4",x"87",x"c7",x"f9"),
   189 => (x"05",x"a8",x"c1",x"86"),
   190 => (x"c2",x"4b",x"87",x"c1"),
   191 => (x"87",x"c5",x"05",x"ab"),
   192 => (x"f9",x"c0",x"48",x"c0"),
   193 => (x"05",x"8b",x"c1",x"87"),
   194 => (x"fc",x"87",x"d0",x"ff"),
   195 => (x"dd",x"c2",x"87",x"f7"),
   196 => (x"98",x"70",x"58",x"ec"),
   197 => (x"c1",x"87",x"cd",x"05"),
   198 => (x"f0",x"ff",x"c0",x"1e"),
   199 => (x"f8",x"49",x"d0",x"c1"),
   200 => (x"86",x"c4",x"87",x"d8"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"de",x"c4",x"78",x"ff"),
   203 => (x"f0",x"dd",x"c2",x"87"),
   204 => (x"48",x"d0",x"ff",x"58"),
   205 => (x"d4",x"ff",x"78",x"c2"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"f5",x"f7",x"48",x"c1"),
   208 => (x"5b",x"5e",x"0e",x"87"),
   209 => (x"71",x"0e",x"5d",x"5c"),
   210 => (x"4d",x"ff",x"c3",x"4a"),
   211 => (x"75",x"4c",x"d4",x"ff"),
   212 => (x"48",x"d0",x"ff",x"7c"),
   213 => (x"75",x"78",x"c3",x"c4"),
   214 => (x"c0",x"1e",x"72",x"7c"),
   215 => (x"d8",x"c1",x"f0",x"ff"),
   216 => (x"87",x"d6",x"f7",x"49"),
   217 => (x"98",x"70",x"86",x"c4"),
   218 => (x"c1",x"87",x"c5",x"02"),
   219 => (x"87",x"f0",x"c0",x"48"),
   220 => (x"fe",x"c3",x"7c",x"75"),
   221 => (x"1e",x"c0",x"c8",x"7c"),
   222 => (x"f4",x"49",x"66",x"d4"),
   223 => (x"86",x"c4",x"87",x"fa"),
   224 => (x"7c",x"75",x"7c",x"75"),
   225 => (x"da",x"d8",x"7c",x"75"),
   226 => (x"7c",x"75",x"4b",x"e0"),
   227 => (x"05",x"99",x"49",x"6c"),
   228 => (x"8b",x"c1",x"87",x"c5"),
   229 => (x"75",x"87",x"f3",x"05"),
   230 => (x"48",x"d0",x"ff",x"7c"),
   231 => (x"48",x"c0",x"78",x"c2"),
   232 => (x"0e",x"87",x"cf",x"f6"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"4b",x"71",x"0e"),
   235 => (x"cd",x"ee",x"c5",x"4c"),
   236 => (x"d4",x"ff",x"4a",x"df"),
   237 => (x"78",x"ff",x"c3",x"48"),
   238 => (x"fe",x"c3",x"49",x"68"),
   239 => (x"fd",x"c0",x"05",x"a9"),
   240 => (x"73",x"4d",x"70",x"87"),
   241 => (x"87",x"cc",x"02",x"9b"),
   242 => (x"73",x"1e",x"66",x"d0"),
   243 => (x"87",x"cf",x"f4",x"49"),
   244 => (x"87",x"d6",x"86",x"c4"),
   245 => (x"c4",x"48",x"d0",x"ff"),
   246 => (x"ff",x"c3",x"78",x"d1"),
   247 => (x"48",x"66",x"d0",x"7d"),
   248 => (x"a6",x"d4",x"88",x"c1"),
   249 => (x"05",x"98",x"70",x"58"),
   250 => (x"d4",x"ff",x"87",x"f0"),
   251 => (x"78",x"ff",x"c3",x"48"),
   252 => (x"05",x"9b",x"73",x"78"),
   253 => (x"d0",x"ff",x"87",x"c5"),
   254 => (x"c1",x"78",x"d0",x"48"),
   255 => (x"8a",x"c1",x"4c",x"4a"),
   256 => (x"87",x"ee",x"fe",x"05"),
   257 => (x"e9",x"f4",x"48",x"74"),
   258 => (x"1e",x"73",x"1e",x"87"),
   259 => (x"4b",x"c0",x"4a",x"71"),
   260 => (x"c3",x"48",x"d4",x"ff"),
   261 => (x"d0",x"ff",x"78",x"ff"),
   262 => (x"78",x"c3",x"c4",x"48"),
   263 => (x"c3",x"48",x"d4",x"ff"),
   264 => (x"1e",x"72",x"78",x"ff"),
   265 => (x"c1",x"f0",x"ff",x"c0"),
   266 => (x"cd",x"f4",x"49",x"d1"),
   267 => (x"70",x"86",x"c4",x"87"),
   268 => (x"87",x"d2",x"05",x"98"),
   269 => (x"cc",x"1e",x"c0",x"c8"),
   270 => (x"e6",x"fd",x"49",x"66"),
   271 => (x"70",x"86",x"c4",x"87"),
   272 => (x"48",x"d0",x"ff",x"4b"),
   273 => (x"48",x"73",x"78",x"c2"),
   274 => (x"0e",x"87",x"eb",x"f3"),
   275 => (x"5d",x"5c",x"5b",x"5e"),
   276 => (x"c0",x"1e",x"c0",x"0e"),
   277 => (x"c9",x"c1",x"f0",x"ff"),
   278 => (x"87",x"de",x"f3",x"49"),
   279 => (x"dd",x"c2",x"1e",x"d2"),
   280 => (x"fe",x"fc",x"49",x"f0"),
   281 => (x"c0",x"86",x"c8",x"87"),
   282 => (x"d2",x"84",x"c1",x"4c"),
   283 => (x"f8",x"04",x"ac",x"b7"),
   284 => (x"f0",x"dd",x"c2",x"87"),
   285 => (x"c3",x"49",x"bf",x"97"),
   286 => (x"c0",x"c1",x"99",x"c0"),
   287 => (x"e7",x"c0",x"05",x"a9"),
   288 => (x"f7",x"dd",x"c2",x"87"),
   289 => (x"d0",x"49",x"bf",x"97"),
   290 => (x"f8",x"dd",x"c2",x"31"),
   291 => (x"c8",x"4a",x"bf",x"97"),
   292 => (x"c2",x"b1",x"72",x"32"),
   293 => (x"bf",x"97",x"f9",x"dd"),
   294 => (x"4c",x"71",x"b1",x"4a"),
   295 => (x"ff",x"ff",x"ff",x"cf"),
   296 => (x"ca",x"84",x"c1",x"9c"),
   297 => (x"87",x"e7",x"c1",x"34"),
   298 => (x"97",x"f9",x"dd",x"c2"),
   299 => (x"31",x"c1",x"49",x"bf"),
   300 => (x"dd",x"c2",x"99",x"c6"),
   301 => (x"4a",x"bf",x"97",x"fa"),
   302 => (x"72",x"2a",x"b7",x"c7"),
   303 => (x"f5",x"dd",x"c2",x"b1"),
   304 => (x"4d",x"4a",x"bf",x"97"),
   305 => (x"dd",x"c2",x"9d",x"cf"),
   306 => (x"4a",x"bf",x"97",x"f6"),
   307 => (x"32",x"ca",x"9a",x"c3"),
   308 => (x"97",x"f7",x"dd",x"c2"),
   309 => (x"33",x"c2",x"4b",x"bf"),
   310 => (x"dd",x"c2",x"b2",x"73"),
   311 => (x"4b",x"bf",x"97",x"f8"),
   312 => (x"c6",x"9b",x"c0",x"c3"),
   313 => (x"b2",x"73",x"2b",x"b7"),
   314 => (x"48",x"c1",x"81",x"c2"),
   315 => (x"49",x"70",x"30",x"71"),
   316 => (x"30",x"75",x"48",x"c1"),
   317 => (x"4c",x"72",x"4d",x"70"),
   318 => (x"94",x"71",x"84",x"c1"),
   319 => (x"ad",x"b7",x"c0",x"c8"),
   320 => (x"c1",x"87",x"cc",x"06"),
   321 => (x"c8",x"2d",x"b7",x"34"),
   322 => (x"01",x"ad",x"b7",x"c0"),
   323 => (x"74",x"87",x"f4",x"ff"),
   324 => (x"87",x"de",x"f0",x"48"),
   325 => (x"5c",x"5b",x"5e",x"0e"),
   326 => (x"86",x"f8",x"0e",x"5d"),
   327 => (x"48",x"d6",x"e6",x"c2"),
   328 => (x"de",x"c2",x"78",x"c0"),
   329 => (x"49",x"c0",x"1e",x"ce"),
   330 => (x"c4",x"87",x"de",x"fb"),
   331 => (x"05",x"98",x"70",x"86"),
   332 => (x"48",x"c0",x"87",x"c5"),
   333 => (x"c0",x"87",x"ce",x"c9"),
   334 => (x"c0",x"7e",x"c1",x"4d"),
   335 => (x"49",x"bf",x"ed",x"f2"),
   336 => (x"4a",x"c4",x"df",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"e0"),
   339 => (x"c0",x"87",x"c2",x"05"),
   340 => (x"e9",x"f2",x"c0",x"7e"),
   341 => (x"df",x"c2",x"49",x"bf"),
   342 => (x"c8",x"71",x"4a",x"e0"),
   343 => (x"87",x"ca",x"ec",x"4b"),
   344 => (x"c2",x"05",x"98",x"70"),
   345 => (x"6e",x"7e",x"c0",x"87"),
   346 => (x"87",x"fd",x"c0",x"02"),
   347 => (x"bf",x"d4",x"e5",x"c2"),
   348 => (x"cc",x"e6",x"c2",x"4d"),
   349 => (x"48",x"7e",x"bf",x"9f"),
   350 => (x"a8",x"ea",x"d6",x"c5"),
   351 => (x"c2",x"87",x"c7",x"05"),
   352 => (x"4d",x"bf",x"d4",x"e5"),
   353 => (x"48",x"6e",x"87",x"ce"),
   354 => (x"a8",x"d5",x"e9",x"ca"),
   355 => (x"c0",x"87",x"c5",x"02"),
   356 => (x"87",x"f1",x"c7",x"48"),
   357 => (x"1e",x"ce",x"de",x"c2"),
   358 => (x"ec",x"f9",x"49",x"75"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"dc",x"c7",x"48",x"c0"),
   362 => (x"e9",x"f2",x"c0",x"87"),
   363 => (x"df",x"c2",x"49",x"bf"),
   364 => (x"c8",x"71",x"4a",x"e0"),
   365 => (x"87",x"f2",x"ea",x"4b"),
   366 => (x"c8",x"05",x"98",x"70"),
   367 => (x"d6",x"e6",x"c2",x"87"),
   368 => (x"da",x"78",x"c1",x"48"),
   369 => (x"ed",x"f2",x"c0",x"87"),
   370 => (x"df",x"c2",x"49",x"bf"),
   371 => (x"c8",x"71",x"4a",x"c4"),
   372 => (x"87",x"d6",x"ea",x"4b"),
   373 => (x"c0",x"02",x"98",x"70"),
   374 => (x"48",x"c0",x"87",x"c5"),
   375 => (x"c2",x"87",x"e6",x"c6"),
   376 => (x"bf",x"97",x"cc",x"e6"),
   377 => (x"a9",x"d5",x"c1",x"49"),
   378 => (x"87",x"cd",x"c0",x"05"),
   379 => (x"97",x"cd",x"e6",x"c2"),
   380 => (x"ea",x"c2",x"49",x"bf"),
   381 => (x"c5",x"c0",x"02",x"a9"),
   382 => (x"c6",x"48",x"c0",x"87"),
   383 => (x"de",x"c2",x"87",x"c7"),
   384 => (x"7e",x"bf",x"97",x"ce"),
   385 => (x"a8",x"e9",x"c3",x"48"),
   386 => (x"87",x"ce",x"c0",x"02"),
   387 => (x"eb",x"c3",x"48",x"6e"),
   388 => (x"c5",x"c0",x"02",x"a8"),
   389 => (x"c5",x"48",x"c0",x"87"),
   390 => (x"de",x"c2",x"87",x"eb"),
   391 => (x"49",x"bf",x"97",x"d9"),
   392 => (x"cc",x"c0",x"05",x"99"),
   393 => (x"da",x"de",x"c2",x"87"),
   394 => (x"c2",x"49",x"bf",x"97"),
   395 => (x"c5",x"c0",x"02",x"a9"),
   396 => (x"c5",x"48",x"c0",x"87"),
   397 => (x"de",x"c2",x"87",x"cf"),
   398 => (x"48",x"bf",x"97",x"db"),
   399 => (x"58",x"d2",x"e6",x"c2"),
   400 => (x"c1",x"48",x"4c",x"70"),
   401 => (x"d6",x"e6",x"c2",x"88"),
   402 => (x"dc",x"de",x"c2",x"58"),
   403 => (x"75",x"49",x"bf",x"97"),
   404 => (x"dd",x"de",x"c2",x"81"),
   405 => (x"c8",x"4a",x"bf",x"97"),
   406 => (x"7e",x"a1",x"72",x"32"),
   407 => (x"48",x"e3",x"ea",x"c2"),
   408 => (x"de",x"c2",x"78",x"6e"),
   409 => (x"48",x"bf",x"97",x"de"),
   410 => (x"c2",x"58",x"a6",x"c8"),
   411 => (x"02",x"bf",x"d6",x"e6"),
   412 => (x"c0",x"87",x"d4",x"c2"),
   413 => (x"49",x"bf",x"e9",x"f2"),
   414 => (x"4a",x"e0",x"df",x"c2"),
   415 => (x"e7",x"4b",x"c8",x"71"),
   416 => (x"98",x"70",x"87",x"e8"),
   417 => (x"87",x"c5",x"c0",x"02"),
   418 => (x"f8",x"c3",x"48",x"c0"),
   419 => (x"ce",x"e6",x"c2",x"87"),
   420 => (x"ea",x"c2",x"4c",x"bf"),
   421 => (x"de",x"c2",x"5c",x"f7"),
   422 => (x"49",x"bf",x"97",x"f3"),
   423 => (x"de",x"c2",x"31",x"c8"),
   424 => (x"4a",x"bf",x"97",x"f2"),
   425 => (x"de",x"c2",x"49",x"a1"),
   426 => (x"4a",x"bf",x"97",x"f4"),
   427 => (x"a1",x"72",x"32",x"d0"),
   428 => (x"f5",x"de",x"c2",x"49"),
   429 => (x"d8",x"4a",x"bf",x"97"),
   430 => (x"49",x"a1",x"72",x"32"),
   431 => (x"c2",x"91",x"66",x"c4"),
   432 => (x"81",x"bf",x"e3",x"ea"),
   433 => (x"59",x"eb",x"ea",x"c2"),
   434 => (x"97",x"fb",x"de",x"c2"),
   435 => (x"32",x"c8",x"4a",x"bf"),
   436 => (x"97",x"fa",x"de",x"c2"),
   437 => (x"4a",x"a2",x"4b",x"bf"),
   438 => (x"97",x"fc",x"de",x"c2"),
   439 => (x"33",x"d0",x"4b",x"bf"),
   440 => (x"c2",x"4a",x"a2",x"73"),
   441 => (x"bf",x"97",x"fd",x"de"),
   442 => (x"d8",x"9b",x"cf",x"4b"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"5a",x"ef",x"ea",x"c2"),
   445 => (x"bf",x"eb",x"ea",x"c2"),
   446 => (x"74",x"8a",x"c2",x"4a"),
   447 => (x"ef",x"ea",x"c2",x"92"),
   448 => (x"78",x"a1",x"72",x"48"),
   449 => (x"c2",x"87",x"ca",x"c1"),
   450 => (x"bf",x"97",x"e0",x"de"),
   451 => (x"c2",x"31",x"c8",x"49"),
   452 => (x"bf",x"97",x"df",x"de"),
   453 => (x"c2",x"49",x"a1",x"4a"),
   454 => (x"c2",x"59",x"de",x"e6"),
   455 => (x"49",x"bf",x"da",x"e6"),
   456 => (x"ff",x"c7",x"31",x"c5"),
   457 => (x"c2",x"29",x"c9",x"81"),
   458 => (x"c2",x"59",x"f7",x"ea"),
   459 => (x"bf",x"97",x"e5",x"de"),
   460 => (x"c2",x"32",x"c8",x"4a"),
   461 => (x"bf",x"97",x"e4",x"de"),
   462 => (x"c4",x"4a",x"a2",x"4b"),
   463 => (x"82",x"6e",x"92",x"66"),
   464 => (x"5a",x"f3",x"ea",x"c2"),
   465 => (x"48",x"eb",x"ea",x"c2"),
   466 => (x"ea",x"c2",x"78",x"c0"),
   467 => (x"a1",x"72",x"48",x"e7"),
   468 => (x"f7",x"ea",x"c2",x"78"),
   469 => (x"eb",x"ea",x"c2",x"48"),
   470 => (x"ea",x"c2",x"78",x"bf"),
   471 => (x"ea",x"c2",x"48",x"fb"),
   472 => (x"c2",x"78",x"bf",x"ef"),
   473 => (x"02",x"bf",x"d6",x"e6"),
   474 => (x"74",x"87",x"c9",x"c0"),
   475 => (x"70",x"30",x"c4",x"48"),
   476 => (x"87",x"c9",x"c0",x"7e"),
   477 => (x"bf",x"f3",x"ea",x"c2"),
   478 => (x"70",x"30",x"c4",x"48"),
   479 => (x"da",x"e6",x"c2",x"7e"),
   480 => (x"c1",x"78",x"6e",x"48"),
   481 => (x"26",x"8e",x"f8",x"48"),
   482 => (x"26",x"4c",x"26",x"4d"),
   483 => (x"0e",x"4f",x"26",x"4b"),
   484 => (x"5d",x"5c",x"5b",x"5e"),
   485 => (x"c2",x"4a",x"71",x"0e"),
   486 => (x"02",x"bf",x"d6",x"e6"),
   487 => (x"4b",x"72",x"87",x"cb"),
   488 => (x"4c",x"72",x"2b",x"c7"),
   489 => (x"c9",x"9c",x"ff",x"c1"),
   490 => (x"c8",x"4b",x"72",x"87"),
   491 => (x"c3",x"4c",x"72",x"2b"),
   492 => (x"ea",x"c2",x"9c",x"ff"),
   493 => (x"c0",x"83",x"bf",x"e3"),
   494 => (x"ab",x"bf",x"e5",x"f2"),
   495 => (x"c0",x"87",x"d9",x"02"),
   496 => (x"c2",x"5b",x"e9",x"f2"),
   497 => (x"73",x"1e",x"ce",x"de"),
   498 => (x"87",x"fd",x"f0",x"49"),
   499 => (x"98",x"70",x"86",x"c4"),
   500 => (x"c0",x"87",x"c5",x"05"),
   501 => (x"87",x"e6",x"c0",x"48"),
   502 => (x"bf",x"d6",x"e6",x"c2"),
   503 => (x"74",x"87",x"d2",x"02"),
   504 => (x"c2",x"91",x"c4",x"49"),
   505 => (x"69",x"81",x"ce",x"de"),
   506 => (x"ff",x"ff",x"cf",x"4d"),
   507 => (x"cb",x"9d",x"ff",x"ff"),
   508 => (x"c2",x"49",x"74",x"87"),
   509 => (x"ce",x"de",x"c2",x"91"),
   510 => (x"4d",x"69",x"9f",x"81"),
   511 => (x"c6",x"fe",x"48",x"75"),
   512 => (x"5b",x"5e",x"0e",x"87"),
   513 => (x"f8",x"0e",x"5d",x"5c"),
   514 => (x"9c",x"4c",x"71",x"86"),
   515 => (x"c0",x"87",x"c5",x"05"),
   516 => (x"87",x"c1",x"c3",x"48"),
   517 => (x"6e",x"7e",x"a4",x"c8"),
   518 => (x"d8",x"78",x"c0",x"48"),
   519 => (x"87",x"c7",x"02",x"66"),
   520 => (x"bf",x"97",x"66",x"d8"),
   521 => (x"c0",x"87",x"c5",x"05"),
   522 => (x"87",x"e9",x"c2",x"48"),
   523 => (x"49",x"c1",x"1e",x"c0"),
   524 => (x"c4",x"87",x"d7",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"de",x"e6",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c9"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ee"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"d5",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"d6",x"e6"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ed"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"d2",x"e6",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fc",x"f9"),
   581 => (x"ce",x"e6",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"d2",x"e6",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d3",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"e7",x"ea",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"ce",x"e6",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"d2",x"e6",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"e9",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d6",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c8",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"e7",x"ea",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"ce",x"e6",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"d2",x"e6",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"e9"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"ff"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f9"),
   629 => (x"0e",x"5d",x"5c",x"5b"),
   630 => (x"d4",x"4b",x"71",x"1e"),
   631 => (x"9b",x"73",x"4d",x"66"),
   632 => (x"87",x"cc",x"c1",x"02"),
   633 => (x"69",x"49",x"a3",x"c8"),
   634 => (x"87",x"c4",x"c1",x"02"),
   635 => (x"c2",x"4c",x"a3",x"d0"),
   636 => (x"49",x"bf",x"d2",x"e6"),
   637 => (x"4a",x"6c",x"b9",x"ff"),
   638 => (x"66",x"d4",x"7e",x"99"),
   639 => (x"87",x"cd",x"06",x"a9"),
   640 => (x"cc",x"7c",x"7b",x"c0"),
   641 => (x"a3",x"c4",x"4a",x"a3"),
   642 => (x"ca",x"79",x"6a",x"49"),
   643 => (x"f8",x"49",x"72",x"87"),
   644 => (x"66",x"d4",x"99",x"c0"),
   645 => (x"75",x"8d",x"71",x"4d"),
   646 => (x"71",x"29",x"c9",x"49"),
   647 => (x"fa",x"49",x"73",x"1e"),
   648 => (x"de",x"c2",x"87",x"f8"),
   649 => (x"49",x"73",x"1e",x"ce"),
   650 => (x"c8",x"87",x"c9",x"fc"),
   651 => (x"7c",x"66",x"d4",x"86"),
   652 => (x"87",x"d3",x"f5",x"26"),
   653 => (x"71",x"1e",x"73",x"1e"),
   654 => (x"c0",x"02",x"9b",x"4b"),
   655 => (x"ea",x"c2",x"87",x"e4"),
   656 => (x"4a",x"73",x"5b",x"fb"),
   657 => (x"e6",x"c2",x"8a",x"c2"),
   658 => (x"92",x"49",x"bf",x"ce"),
   659 => (x"bf",x"e7",x"ea",x"c2"),
   660 => (x"c2",x"80",x"72",x"48"),
   661 => (x"71",x"58",x"ff",x"ea"),
   662 => (x"c2",x"30",x"c4",x"48"),
   663 => (x"c0",x"58",x"de",x"e6"),
   664 => (x"ea",x"c2",x"87",x"ed"),
   665 => (x"ea",x"c2",x"48",x"f7"),
   666 => (x"c2",x"78",x"bf",x"eb"),
   667 => (x"c2",x"48",x"fb",x"ea"),
   668 => (x"78",x"bf",x"ef",x"ea"),
   669 => (x"bf",x"d6",x"e6",x"c2"),
   670 => (x"c2",x"87",x"c9",x"02"),
   671 => (x"49",x"bf",x"ce",x"e6"),
   672 => (x"87",x"c7",x"31",x"c4"),
   673 => (x"bf",x"f3",x"ea",x"c2"),
   674 => (x"c2",x"31",x"c4",x"49"),
   675 => (x"f3",x"59",x"de",x"e6"),
   676 => (x"5e",x"0e",x"87",x"f9"),
   677 => (x"71",x"0e",x"5c",x"5b"),
   678 => (x"72",x"4b",x"c0",x"4a"),
   679 => (x"e1",x"c0",x"02",x"9a"),
   680 => (x"49",x"a2",x"da",x"87"),
   681 => (x"c2",x"4b",x"69",x"9f"),
   682 => (x"02",x"bf",x"d6",x"e6"),
   683 => (x"a2",x"d4",x"87",x"cf"),
   684 => (x"49",x"69",x"9f",x"49"),
   685 => (x"ff",x"ff",x"c0",x"4c"),
   686 => (x"c2",x"34",x"d0",x"9c"),
   687 => (x"74",x"4c",x"c0",x"87"),
   688 => (x"49",x"73",x"b3",x"49"),
   689 => (x"f2",x"87",x"ed",x"fd"),
   690 => (x"5e",x"0e",x"87",x"ff"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4a",x"71",x"86",x"f4"),
   693 => (x"9a",x"72",x"7e",x"c0"),
   694 => (x"c2",x"87",x"d8",x"02"),
   695 => (x"c0",x"48",x"ca",x"de"),
   696 => (x"c2",x"de",x"c2",x"78"),
   697 => (x"fb",x"ea",x"c2",x"48"),
   698 => (x"de",x"c2",x"78",x"bf"),
   699 => (x"ea",x"c2",x"48",x"c6"),
   700 => (x"c2",x"78",x"bf",x"f7"),
   701 => (x"c0",x"48",x"eb",x"e6"),
   702 => (x"da",x"e6",x"c2",x"50"),
   703 => (x"de",x"c2",x"49",x"bf"),
   704 => (x"71",x"4a",x"bf",x"ca"),
   705 => (x"c9",x"c4",x"03",x"aa"),
   706 => (x"cf",x"49",x"72",x"87"),
   707 => (x"e9",x"c0",x"05",x"99"),
   708 => (x"e5",x"f2",x"c0",x"87"),
   709 => (x"c2",x"de",x"c2",x"48"),
   710 => (x"de",x"c2",x"78",x"bf"),
   711 => (x"de",x"c2",x"1e",x"ce"),
   712 => (x"c2",x"49",x"bf",x"c2"),
   713 => (x"c1",x"48",x"c2",x"de"),
   714 => (x"e3",x"71",x"78",x"a1"),
   715 => (x"86",x"c4",x"87",x"db"),
   716 => (x"48",x"e1",x"f2",x"c0"),
   717 => (x"78",x"ce",x"de",x"c2"),
   718 => (x"f2",x"c0",x"87",x"cc"),
   719 => (x"c0",x"48",x"bf",x"e1"),
   720 => (x"f2",x"c0",x"80",x"e0"),
   721 => (x"de",x"c2",x"58",x"e5"),
   722 => (x"c1",x"48",x"bf",x"ca"),
   723 => (x"ce",x"de",x"c2",x"80"),
   724 => (x"0c",x"a1",x"27",x"58"),
   725 => (x"97",x"bf",x"00",x"00"),
   726 => (x"02",x"9d",x"4d",x"bf"),
   727 => (x"c3",x"87",x"e3",x"c2"),
   728 => (x"c2",x"02",x"ad",x"e5"),
   729 => (x"f2",x"c0",x"87",x"dc"),
   730 => (x"cb",x"4b",x"bf",x"e1"),
   731 => (x"4c",x"11",x"49",x"a3"),
   732 => (x"c1",x"05",x"ac",x"cf"),
   733 => (x"49",x"75",x"87",x"d2"),
   734 => (x"89",x"c1",x"99",x"df"),
   735 => (x"e6",x"c2",x"91",x"cd"),
   736 => (x"a3",x"c1",x"81",x"de"),
   737 => (x"c3",x"51",x"12",x"4a"),
   738 => (x"51",x"12",x"4a",x"a3"),
   739 => (x"12",x"4a",x"a3",x"c5"),
   740 => (x"4a",x"a3",x"c7",x"51"),
   741 => (x"a3",x"c9",x"51",x"12"),
   742 => (x"ce",x"51",x"12",x"4a"),
   743 => (x"51",x"12",x"4a",x"a3"),
   744 => (x"12",x"4a",x"a3",x"d0"),
   745 => (x"4a",x"a3",x"d2",x"51"),
   746 => (x"a3",x"d4",x"51",x"12"),
   747 => (x"d6",x"51",x"12",x"4a"),
   748 => (x"51",x"12",x"4a",x"a3"),
   749 => (x"12",x"4a",x"a3",x"d8"),
   750 => (x"4a",x"a3",x"dc",x"51"),
   751 => (x"a3",x"de",x"51",x"12"),
   752 => (x"c1",x"51",x"12",x"4a"),
   753 => (x"87",x"fa",x"c0",x"7e"),
   754 => (x"99",x"c8",x"49",x"74"),
   755 => (x"87",x"eb",x"c0",x"05"),
   756 => (x"99",x"d0",x"49",x"74"),
   757 => (x"dc",x"87",x"d1",x"05"),
   758 => (x"cb",x"c0",x"02",x"66"),
   759 => (x"dc",x"49",x"73",x"87"),
   760 => (x"98",x"70",x"0f",x"66"),
   761 => (x"87",x"d3",x"c0",x"02"),
   762 => (x"c6",x"c0",x"05",x"6e"),
   763 => (x"de",x"e6",x"c2",x"87"),
   764 => (x"c0",x"50",x"c0",x"48"),
   765 => (x"48",x"bf",x"e1",x"f2"),
   766 => (x"c2",x"87",x"e1",x"c2"),
   767 => (x"c0",x"48",x"eb",x"e6"),
   768 => (x"e6",x"c2",x"7e",x"50"),
   769 => (x"c2",x"49",x"bf",x"da"),
   770 => (x"4a",x"bf",x"ca",x"de"),
   771 => (x"fb",x"04",x"aa",x"71"),
   772 => (x"ea",x"c2",x"87",x"f7"),
   773 => (x"c0",x"05",x"bf",x"fb"),
   774 => (x"e6",x"c2",x"87",x"c8"),
   775 => (x"c1",x"02",x"bf",x"d6"),
   776 => (x"de",x"c2",x"87",x"f8"),
   777 => (x"ed",x"49",x"bf",x"c6"),
   778 => (x"49",x"70",x"87",x"e5"),
   779 => (x"59",x"ca",x"de",x"c2"),
   780 => (x"c2",x"48",x"a6",x"c4"),
   781 => (x"78",x"bf",x"c6",x"de"),
   782 => (x"bf",x"d6",x"e6",x"c2"),
   783 => (x"87",x"d8",x"c0",x"02"),
   784 => (x"cf",x"49",x"66",x"c4"),
   785 => (x"f8",x"ff",x"ff",x"ff"),
   786 => (x"c0",x"02",x"a9",x"99"),
   787 => (x"4c",x"c0",x"87",x"c5"),
   788 => (x"c1",x"87",x"e1",x"c0"),
   789 => (x"87",x"dc",x"c0",x"4c"),
   790 => (x"cf",x"49",x"66",x"c4"),
   791 => (x"a9",x"99",x"f8",x"ff"),
   792 => (x"87",x"c8",x"c0",x"02"),
   793 => (x"c0",x"48",x"a6",x"c8"),
   794 => (x"87",x"c5",x"c0",x"78"),
   795 => (x"c1",x"48",x"a6",x"c8"),
   796 => (x"4c",x"66",x"c8",x"78"),
   797 => (x"c0",x"05",x"9c",x"74"),
   798 => (x"66",x"c4",x"87",x"e0"),
   799 => (x"c2",x"89",x"c2",x"49"),
   800 => (x"4a",x"bf",x"ce",x"e6"),
   801 => (x"e7",x"ea",x"c2",x"91"),
   802 => (x"de",x"c2",x"4a",x"bf"),
   803 => (x"a1",x"72",x"48",x"c2"),
   804 => (x"ca",x"de",x"c2",x"78"),
   805 => (x"f9",x"78",x"c0",x"48"),
   806 => (x"48",x"c0",x"87",x"df"),
   807 => (x"e6",x"eb",x"8e",x"f4"),
   808 => (x"00",x"00",x"00",x"87"),
   809 => (x"ff",x"ff",x"ff",x"00"),
   810 => (x"00",x"0c",x"b1",x"ff"),
   811 => (x"00",x"0c",x"ba",x"00"),
   812 => (x"54",x"41",x"46",x"00"),
   813 => (x"20",x"20",x"32",x"33"),
   814 => (x"41",x"46",x"00",x"20"),
   815 => (x"20",x"36",x"31",x"54"),
   816 => (x"1e",x"00",x"20",x"20"),
   817 => (x"c3",x"48",x"d4",x"ff"),
   818 => (x"48",x"68",x"78",x"ff"),
   819 => (x"ff",x"1e",x"4f",x"26"),
   820 => (x"ff",x"c3",x"48",x"d4"),
   821 => (x"48",x"d0",x"ff",x"78"),
   822 => (x"ff",x"78",x"e1",x"c0"),
   823 => (x"78",x"d4",x"48",x"d4"),
   824 => (x"48",x"ff",x"ea",x"c2"),
   825 => (x"50",x"bf",x"d4",x"ff"),
   826 => (x"ff",x"1e",x"4f",x"26"),
   827 => (x"e0",x"c0",x"48",x"d0"),
   828 => (x"1e",x"4f",x"26",x"78"),
   829 => (x"70",x"87",x"cc",x"ff"),
   830 => (x"c6",x"02",x"99",x"49"),
   831 => (x"a9",x"fb",x"c0",x"87"),
   832 => (x"71",x"87",x"f1",x"05"),
   833 => (x"0e",x"4f",x"26",x"48"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"4c",x"c0",x"4b",x"71"),
   836 => (x"70",x"87",x"f0",x"fe"),
   837 => (x"c0",x"02",x"99",x"49"),
   838 => (x"ec",x"c0",x"87",x"f9"),
   839 => (x"f2",x"c0",x"02",x"a9"),
   840 => (x"a9",x"fb",x"c0",x"87"),
   841 => (x"87",x"eb",x"c0",x"02"),
   842 => (x"ac",x"b7",x"66",x"cc"),
   843 => (x"d0",x"87",x"c7",x"03"),
   844 => (x"87",x"c2",x"02",x"66"),
   845 => (x"99",x"71",x"53",x"71"),
   846 => (x"c1",x"87",x"c2",x"02"),
   847 => (x"87",x"c3",x"fe",x"84"),
   848 => (x"02",x"99",x"49",x"70"),
   849 => (x"ec",x"c0",x"87",x"cd"),
   850 => (x"87",x"c7",x"02",x"a9"),
   851 => (x"05",x"a9",x"fb",x"c0"),
   852 => (x"d0",x"87",x"d5",x"ff"),
   853 => (x"87",x"c3",x"02",x"66"),
   854 => (x"c0",x"7b",x"97",x"c0"),
   855 => (x"c4",x"05",x"a9",x"ec"),
   856 => (x"c5",x"4a",x"74",x"87"),
   857 => (x"c0",x"4a",x"74",x"87"),
   858 => (x"48",x"72",x"8a",x"0a"),
   859 => (x"4d",x"26",x"87",x"c2"),
   860 => (x"4b",x"26",x"4c",x"26"),
   861 => (x"fd",x"1e",x"4f",x"26"),
   862 => (x"49",x"70",x"87",x"c9"),
   863 => (x"aa",x"f0",x"c0",x"4a"),
   864 => (x"c0",x"87",x"c9",x"04"),
   865 => (x"c3",x"01",x"aa",x"f9"),
   866 => (x"8a",x"f0",x"c0",x"87"),
   867 => (x"04",x"aa",x"c1",x"c1"),
   868 => (x"da",x"c1",x"87",x"c9"),
   869 => (x"87",x"c3",x"01",x"aa"),
   870 => (x"72",x"8a",x"f7",x"c0"),
   871 => (x"0e",x"4f",x"26",x"48"),
   872 => (x"0e",x"5c",x"5b",x"5e"),
   873 => (x"d4",x"ff",x"4a",x"71"),
   874 => (x"c0",x"49",x"72",x"4c"),
   875 => (x"4b",x"70",x"87",x"e9"),
   876 => (x"87",x"c2",x"02",x"9b"),
   877 => (x"d0",x"ff",x"8b",x"c1"),
   878 => (x"c1",x"78",x"c5",x"48"),
   879 => (x"49",x"73",x"7c",x"d5"),
   880 => (x"e3",x"c1",x"31",x"c6"),
   881 => (x"4a",x"bf",x"97",x"d0"),
   882 => (x"70",x"b0",x"71",x"48"),
   883 => (x"48",x"d0",x"ff",x"7c"),
   884 => (x"48",x"73",x"78",x"c4"),
   885 => (x"0e",x"87",x"d9",x"fe"),
   886 => (x"5d",x"5c",x"5b",x"5e"),
   887 => (x"71",x"86",x"f8",x"0e"),
   888 => (x"fb",x"7e",x"c0",x"4c"),
   889 => (x"4b",x"c0",x"87",x"e8"),
   890 => (x"97",x"c4",x"fa",x"c0"),
   891 => (x"a9",x"c0",x"49",x"bf"),
   892 => (x"fb",x"87",x"cf",x"04"),
   893 => (x"83",x"c1",x"87",x"fd"),
   894 => (x"97",x"c4",x"fa",x"c0"),
   895 => (x"06",x"ab",x"49",x"bf"),
   896 => (x"fa",x"c0",x"87",x"f1"),
   897 => (x"02",x"bf",x"97",x"c4"),
   898 => (x"f6",x"fa",x"87",x"cf"),
   899 => (x"99",x"49",x"70",x"87"),
   900 => (x"c0",x"87",x"c6",x"02"),
   901 => (x"f1",x"05",x"a9",x"ec"),
   902 => (x"fa",x"4b",x"c0",x"87"),
   903 => (x"4d",x"70",x"87",x"e5"),
   904 => (x"c8",x"87",x"e0",x"fa"),
   905 => (x"da",x"fa",x"58",x"a6"),
   906 => (x"c1",x"4a",x"70",x"87"),
   907 => (x"49",x"a4",x"c8",x"83"),
   908 => (x"ad",x"49",x"69",x"97"),
   909 => (x"c0",x"87",x"c7",x"02"),
   910 => (x"c0",x"05",x"ad",x"ff"),
   911 => (x"a4",x"c9",x"87",x"e7"),
   912 => (x"49",x"69",x"97",x"49"),
   913 => (x"02",x"a9",x"66",x"c4"),
   914 => (x"c0",x"48",x"87",x"c7"),
   915 => (x"d4",x"05",x"a8",x"ff"),
   916 => (x"49",x"a4",x"ca",x"87"),
   917 => (x"aa",x"49",x"69",x"97"),
   918 => (x"c0",x"87",x"c6",x"02"),
   919 => (x"c4",x"05",x"aa",x"ff"),
   920 => (x"d0",x"7e",x"c1",x"87"),
   921 => (x"ad",x"ec",x"c0",x"87"),
   922 => (x"c0",x"87",x"c6",x"02"),
   923 => (x"c4",x"05",x"ad",x"fb"),
   924 => (x"c1",x"4b",x"c0",x"87"),
   925 => (x"fe",x"02",x"6e",x"7e"),
   926 => (x"ed",x"f9",x"87",x"e1"),
   927 => (x"f8",x"48",x"73",x"87"),
   928 => (x"87",x"ea",x"fb",x"8e"),
   929 => (x"5b",x"5e",x"0e",x"00"),
   930 => (x"f8",x"0e",x"5d",x"5c"),
   931 => (x"ff",x"4d",x"71",x"86"),
   932 => (x"1e",x"75",x"4b",x"d4"),
   933 => (x"49",x"c4",x"eb",x"c2"),
   934 => (x"c4",x"87",x"e6",x"e5"),
   935 => (x"02",x"98",x"70",x"86"),
   936 => (x"c4",x"87",x"cc",x"c4"),
   937 => (x"e3",x"c1",x"48",x"a6"),
   938 => (x"75",x"78",x"bf",x"d2"),
   939 => (x"87",x"ef",x"fb",x"49"),
   940 => (x"c5",x"48",x"d0",x"ff"),
   941 => (x"7b",x"d6",x"c1",x"78"),
   942 => (x"a2",x"75",x"4a",x"c0"),
   943 => (x"c1",x"7b",x"11",x"49"),
   944 => (x"aa",x"b7",x"cb",x"82"),
   945 => (x"cc",x"87",x"f3",x"04"),
   946 => (x"7b",x"ff",x"c3",x"4a"),
   947 => (x"e0",x"c0",x"82",x"c1"),
   948 => (x"f4",x"04",x"aa",x"b7"),
   949 => (x"48",x"d0",x"ff",x"87"),
   950 => (x"ff",x"c3",x"78",x"c4"),
   951 => (x"c1",x"78",x"c5",x"7b"),
   952 => (x"7b",x"c1",x"7b",x"d3"),
   953 => (x"48",x"66",x"78",x"c4"),
   954 => (x"06",x"a8",x"b7",x"c0"),
   955 => (x"c2",x"87",x"f0",x"c2"),
   956 => (x"4c",x"bf",x"cc",x"eb"),
   957 => (x"74",x"48",x"66",x"c4"),
   958 => (x"58",x"a6",x"c8",x"88"),
   959 => (x"c1",x"02",x"9c",x"74"),
   960 => (x"de",x"c2",x"87",x"f9"),
   961 => (x"c0",x"c8",x"7e",x"ce"),
   962 => (x"b7",x"c0",x"8c",x"4d"),
   963 => (x"87",x"c6",x"03",x"ac"),
   964 => (x"4d",x"a4",x"c0",x"c8"),
   965 => (x"ea",x"c2",x"4c",x"c0"),
   966 => (x"49",x"bf",x"97",x"ff"),
   967 => (x"d1",x"02",x"99",x"d0"),
   968 => (x"c2",x"1e",x"c0",x"87"),
   969 => (x"e8",x"49",x"c4",x"eb"),
   970 => (x"86",x"c4",x"87",x"ca"),
   971 => (x"c0",x"4a",x"49",x"70"),
   972 => (x"de",x"c2",x"87",x"ee"),
   973 => (x"eb",x"c2",x"1e",x"ce"),
   974 => (x"f7",x"e7",x"49",x"c4"),
   975 => (x"70",x"86",x"c4",x"87"),
   976 => (x"d0",x"ff",x"4a",x"49"),
   977 => (x"78",x"c5",x"c8",x"48"),
   978 => (x"6e",x"7b",x"d4",x"c1"),
   979 => (x"6e",x"7b",x"bf",x"97"),
   980 => (x"70",x"80",x"c1",x"48"),
   981 => (x"05",x"8d",x"c1",x"7e"),
   982 => (x"ff",x"87",x"f0",x"ff"),
   983 => (x"78",x"c4",x"48",x"d0"),
   984 => (x"c5",x"05",x"9a",x"72"),
   985 => (x"c1",x"48",x"c0",x"87"),
   986 => (x"1e",x"c1",x"87",x"c7"),
   987 => (x"49",x"c4",x"eb",x"c2"),
   988 => (x"c4",x"87",x"e7",x"e5"),
   989 => (x"05",x"9c",x"74",x"86"),
   990 => (x"c4",x"87",x"c7",x"fe"),
   991 => (x"b7",x"c0",x"48",x"66"),
   992 => (x"87",x"d1",x"06",x"a8"),
   993 => (x"48",x"c4",x"eb",x"c2"),
   994 => (x"80",x"d0",x"78",x"c0"),
   995 => (x"80",x"f4",x"78",x"c0"),
   996 => (x"bf",x"d0",x"eb",x"c2"),
   997 => (x"48",x"66",x"c4",x"78"),
   998 => (x"01",x"a8",x"b7",x"c0"),
   999 => (x"ff",x"87",x"d0",x"fd"),
  1000 => (x"78",x"c5",x"48",x"d0"),
  1001 => (x"c0",x"7b",x"d3",x"c1"),
  1002 => (x"c1",x"78",x"c4",x"7b"),
  1003 => (x"c0",x"87",x"c2",x"48"),
  1004 => (x"26",x"8e",x"f8",x"48"),
  1005 => (x"26",x"4c",x"26",x"4d"),
  1006 => (x"0e",x"4f",x"26",x"4b"),
  1007 => (x"5d",x"5c",x"5b",x"5e"),
  1008 => (x"4b",x"71",x"1e",x"0e"),
  1009 => (x"ab",x"4d",x"4c",x"c0"),
  1010 => (x"87",x"e8",x"c0",x"04"),
  1011 => (x"1e",x"d7",x"f7",x"c0"),
  1012 => (x"c4",x"02",x"9d",x"75"),
  1013 => (x"c2",x"4a",x"c0",x"87"),
  1014 => (x"72",x"4a",x"c1",x"87"),
  1015 => (x"87",x"ea",x"eb",x"49"),
  1016 => (x"7e",x"70",x"86",x"c4"),
  1017 => (x"05",x"6e",x"84",x"c1"),
  1018 => (x"4c",x"73",x"87",x"c2"),
  1019 => (x"ac",x"73",x"85",x"c1"),
  1020 => (x"87",x"d8",x"ff",x"06"),
  1021 => (x"fe",x"26",x"48",x"6e"),
  1022 => (x"5e",x"0e",x"87",x"f9"),
  1023 => (x"71",x"0e",x"5c",x"5b"),
  1024 => (x"02",x"66",x"cc",x"4b"),
  1025 => (x"c0",x"4c",x"87",x"d8"),
  1026 => (x"d8",x"02",x"8c",x"f0"),
  1027 => (x"c1",x"4a",x"74",x"87"),
  1028 => (x"87",x"d1",x"02",x"8a"),
  1029 => (x"87",x"cd",x"02",x"8a"),
  1030 => (x"87",x"c9",x"02",x"8a"),
  1031 => (x"49",x"73",x"87",x"d9"),
  1032 => (x"d2",x"87",x"e2",x"f9"),
  1033 => (x"c0",x"1e",x"74",x"87"),
  1034 => (x"ef",x"d7",x"c1",x"49"),
  1035 => (x"73",x"1e",x"74",x"87"),
  1036 => (x"e7",x"d7",x"c1",x"49"),
  1037 => (x"fd",x"86",x"c8",x"87"),
  1038 => (x"5e",x"0e",x"87",x"fb"),
  1039 => (x"0e",x"5d",x"5c",x"5b"),
  1040 => (x"49",x"4c",x"71",x"1e"),
  1041 => (x"eb",x"c2",x"91",x"de"),
  1042 => (x"85",x"71",x"4d",x"ec"),
  1043 => (x"c1",x"02",x"6d",x"97"),
  1044 => (x"eb",x"c2",x"87",x"dc"),
  1045 => (x"74",x"4a",x"bf",x"d8"),
  1046 => (x"fd",x"49",x"72",x"82"),
  1047 => (x"7e",x"70",x"87",x"dd"),
  1048 => (x"f2",x"c0",x"02",x"6e"),
  1049 => (x"e0",x"eb",x"c2",x"87"),
  1050 => (x"cb",x"4a",x"6e",x"4b"),
  1051 => (x"f7",x"c0",x"ff",x"49"),
  1052 => (x"cb",x"4b",x"74",x"87"),
  1053 => (x"e4",x"e3",x"c1",x"93"),
  1054 => (x"c1",x"83",x"c4",x"83"),
  1055 => (x"74",x"7b",x"f2",x"c2"),
  1056 => (x"f0",x"c1",x"c1",x"49"),
  1057 => (x"c1",x"7b",x"75",x"87"),
  1058 => (x"bf",x"97",x"d1",x"e3"),
  1059 => (x"eb",x"c2",x"1e",x"49"),
  1060 => (x"e5",x"fd",x"49",x"e0"),
  1061 => (x"74",x"86",x"c4",x"87"),
  1062 => (x"d8",x"c1",x"c1",x"49"),
  1063 => (x"c1",x"49",x"c0",x"87"),
  1064 => (x"c2",x"87",x"f7",x"c2"),
  1065 => (x"c0",x"48",x"c0",x"eb"),
  1066 => (x"dd",x"49",x"c1",x"78"),
  1067 => (x"fc",x"26",x"87",x"da"),
  1068 => (x"6f",x"4c",x"87",x"c1"),
  1069 => (x"6e",x"69",x"64",x"61"),
  1070 => (x"2e",x"2e",x"2e",x"67"),
  1071 => (x"5b",x"5e",x"0e",x"00"),
  1072 => (x"4b",x"71",x"0e",x"5c"),
  1073 => (x"d8",x"eb",x"c2",x"4a"),
  1074 => (x"49",x"72",x"82",x"bf"),
  1075 => (x"70",x"87",x"ec",x"fb"),
  1076 => (x"c4",x"02",x"9c",x"4c"),
  1077 => (x"f9",x"e6",x"49",x"87"),
  1078 => (x"d8",x"eb",x"c2",x"87"),
  1079 => (x"c1",x"78",x"c0",x"48"),
  1080 => (x"87",x"e4",x"dc",x"49"),
  1081 => (x"0e",x"87",x"ce",x"fb"),
  1082 => (x"5d",x"5c",x"5b",x"5e"),
  1083 => (x"c2",x"86",x"f4",x"0e"),
  1084 => (x"c0",x"4d",x"ce",x"de"),
  1085 => (x"48",x"a6",x"c4",x"4c"),
  1086 => (x"eb",x"c2",x"78",x"c0"),
  1087 => (x"c0",x"49",x"bf",x"d8"),
  1088 => (x"c1",x"c1",x"06",x"a9"),
  1089 => (x"ce",x"de",x"c2",x"87"),
  1090 => (x"c0",x"02",x"98",x"48"),
  1091 => (x"f7",x"c0",x"87",x"f8"),
  1092 => (x"66",x"c8",x"1e",x"d7"),
  1093 => (x"c4",x"87",x"c7",x"02"),
  1094 => (x"78",x"c0",x"48",x"a6"),
  1095 => (x"a6",x"c4",x"87",x"c5"),
  1096 => (x"c4",x"78",x"c1",x"48"),
  1097 => (x"e1",x"e6",x"49",x"66"),
  1098 => (x"70",x"86",x"c4",x"87"),
  1099 => (x"c4",x"84",x"c1",x"4d"),
  1100 => (x"80",x"c1",x"48",x"66"),
  1101 => (x"c2",x"58",x"a6",x"c8"),
  1102 => (x"49",x"bf",x"d8",x"eb"),
  1103 => (x"87",x"c6",x"03",x"ac"),
  1104 => (x"ff",x"05",x"9d",x"75"),
  1105 => (x"4c",x"c0",x"87",x"c8"),
  1106 => (x"c3",x"02",x"9d",x"75"),
  1107 => (x"f7",x"c0",x"87",x"e0"),
  1108 => (x"66",x"c8",x"1e",x"d7"),
  1109 => (x"cc",x"87",x"c7",x"02"),
  1110 => (x"78",x"c0",x"48",x"a6"),
  1111 => (x"a6",x"cc",x"87",x"c5"),
  1112 => (x"cc",x"78",x"c1",x"48"),
  1113 => (x"e1",x"e5",x"49",x"66"),
  1114 => (x"70",x"86",x"c4",x"87"),
  1115 => (x"c2",x"02",x"6e",x"7e"),
  1116 => (x"49",x"6e",x"87",x"e9"),
  1117 => (x"69",x"97",x"81",x"cb"),
  1118 => (x"02",x"99",x"d0",x"49"),
  1119 => (x"c1",x"87",x"d6",x"c1"),
  1120 => (x"74",x"4a",x"fd",x"c2"),
  1121 => (x"c1",x"91",x"cb",x"49"),
  1122 => (x"72",x"81",x"e4",x"e3"),
  1123 => (x"c3",x"81",x"c8",x"79"),
  1124 => (x"49",x"74",x"51",x"ff"),
  1125 => (x"eb",x"c2",x"91",x"de"),
  1126 => (x"85",x"71",x"4d",x"ec"),
  1127 => (x"7d",x"97",x"c1",x"c2"),
  1128 => (x"c0",x"49",x"a5",x"c1"),
  1129 => (x"e6",x"c2",x"51",x"e0"),
  1130 => (x"02",x"bf",x"97",x"de"),
  1131 => (x"84",x"c1",x"87",x"d2"),
  1132 => (x"c2",x"4b",x"a5",x"c2"),
  1133 => (x"db",x"4a",x"de",x"e6"),
  1134 => (x"eb",x"fb",x"fe",x"49"),
  1135 => (x"87",x"db",x"c1",x"87"),
  1136 => (x"c0",x"49",x"a5",x"cd"),
  1137 => (x"c2",x"84",x"c1",x"51"),
  1138 => (x"4a",x"6e",x"4b",x"a5"),
  1139 => (x"fb",x"fe",x"49",x"cb"),
  1140 => (x"c6",x"c1",x"87",x"d6"),
  1141 => (x"fa",x"c0",x"c1",x"87"),
  1142 => (x"cb",x"49",x"74",x"4a"),
  1143 => (x"e4",x"e3",x"c1",x"91"),
  1144 => (x"c2",x"79",x"72",x"81"),
  1145 => (x"bf",x"97",x"de",x"e6"),
  1146 => (x"74",x"87",x"d8",x"02"),
  1147 => (x"c1",x"91",x"de",x"49"),
  1148 => (x"ec",x"eb",x"c2",x"84"),
  1149 => (x"c2",x"83",x"71",x"4b"),
  1150 => (x"dd",x"4a",x"de",x"e6"),
  1151 => (x"e7",x"fa",x"fe",x"49"),
  1152 => (x"74",x"87",x"d8",x"87"),
  1153 => (x"c2",x"93",x"de",x"4b"),
  1154 => (x"cb",x"83",x"ec",x"eb"),
  1155 => (x"51",x"c0",x"49",x"a3"),
  1156 => (x"6e",x"73",x"84",x"c1"),
  1157 => (x"fe",x"49",x"cb",x"4a"),
  1158 => (x"c4",x"87",x"cd",x"fa"),
  1159 => (x"80",x"c1",x"48",x"66"),
  1160 => (x"c7",x"58",x"a6",x"c8"),
  1161 => (x"c5",x"c0",x"03",x"ac"),
  1162 => (x"fc",x"05",x"6e",x"87"),
  1163 => (x"48",x"74",x"87",x"e0"),
  1164 => (x"fe",x"f5",x"8e",x"f4"),
  1165 => (x"1e",x"73",x"1e",x"87"),
  1166 => (x"cb",x"49",x"4b",x"71"),
  1167 => (x"e4",x"e3",x"c1",x"91"),
  1168 => (x"4a",x"a1",x"c8",x"81"),
  1169 => (x"48",x"d0",x"e3",x"c1"),
  1170 => (x"a1",x"c9",x"50",x"12"),
  1171 => (x"c4",x"fa",x"c0",x"4a"),
  1172 => (x"ca",x"50",x"12",x"48"),
  1173 => (x"d1",x"e3",x"c1",x"81"),
  1174 => (x"c1",x"50",x"11",x"48"),
  1175 => (x"bf",x"97",x"d1",x"e3"),
  1176 => (x"49",x"c0",x"1e",x"49"),
  1177 => (x"c2",x"87",x"d3",x"f6"),
  1178 => (x"de",x"48",x"c0",x"eb"),
  1179 => (x"d6",x"49",x"c1",x"78"),
  1180 => (x"f5",x"26",x"87",x"d6"),
  1181 => (x"71",x"1e",x"87",x"c1"),
  1182 => (x"91",x"cb",x"49",x"4a"),
  1183 => (x"81",x"e4",x"e3",x"c1"),
  1184 => (x"48",x"11",x"81",x"c8"),
  1185 => (x"58",x"c4",x"eb",x"c2"),
  1186 => (x"48",x"d8",x"eb",x"c2"),
  1187 => (x"49",x"c1",x"78",x"c0"),
  1188 => (x"26",x"87",x"f5",x"d5"),
  1189 => (x"49",x"c0",x"1e",x"4f"),
  1190 => (x"87",x"fe",x"fa",x"c0"),
  1191 => (x"71",x"1e",x"4f",x"26"),
  1192 => (x"87",x"d2",x"02",x"99"),
  1193 => (x"48",x"f9",x"e4",x"c1"),
  1194 => (x"80",x"f7",x"50",x"c0"),
  1195 => (x"40",x"f6",x"c9",x"c1"),
  1196 => (x"78",x"dd",x"e3",x"c1"),
  1197 => (x"e4",x"c1",x"87",x"ce"),
  1198 => (x"e3",x"c1",x"48",x"f5"),
  1199 => (x"80",x"fc",x"78",x"d6"),
  1200 => (x"78",x"d5",x"ca",x"c1"),
  1201 => (x"5e",x"0e",x"4f",x"26"),
  1202 => (x"71",x"0e",x"5c",x"5b"),
  1203 => (x"92",x"cb",x"4a",x"4c"),
  1204 => (x"82",x"e4",x"e3",x"c1"),
  1205 => (x"c9",x"49",x"a2",x"c8"),
  1206 => (x"6b",x"97",x"4b",x"a2"),
  1207 => (x"69",x"97",x"1e",x"4b"),
  1208 => (x"82",x"ca",x"1e",x"49"),
  1209 => (x"e5",x"c0",x"49",x"12"),
  1210 => (x"49",x"c0",x"87",x"f9"),
  1211 => (x"74",x"87",x"d9",x"d4"),
  1212 => (x"c0",x"f8",x"c0",x"49"),
  1213 => (x"f2",x"8e",x"f8",x"87"),
  1214 => (x"73",x"1e",x"87",x"fb"),
  1215 => (x"49",x"4b",x"71",x"1e"),
  1216 => (x"73",x"87",x"c3",x"ff"),
  1217 => (x"87",x"fe",x"fe",x"49"),
  1218 => (x"1e",x"87",x"ec",x"f2"),
  1219 => (x"4b",x"71",x"1e",x"73"),
  1220 => (x"02",x"4a",x"a3",x"c6"),
  1221 => (x"8a",x"c1",x"87",x"db"),
  1222 => (x"8a",x"87",x"d6",x"02"),
  1223 => (x"87",x"da",x"c1",x"02"),
  1224 => (x"fc",x"c0",x"02",x"8a"),
  1225 => (x"c0",x"02",x"8a",x"87"),
  1226 => (x"02",x"8a",x"87",x"e1"),
  1227 => (x"db",x"c1",x"87",x"cb"),
  1228 => (x"fd",x"49",x"c7",x"87"),
  1229 => (x"de",x"c1",x"87",x"c0"),
  1230 => (x"d8",x"eb",x"c2",x"87"),
  1231 => (x"cb",x"c1",x"02",x"bf"),
  1232 => (x"88",x"c1",x"48",x"87"),
  1233 => (x"58",x"dc",x"eb",x"c2"),
  1234 => (x"c2",x"87",x"c1",x"c1"),
  1235 => (x"02",x"bf",x"dc",x"eb"),
  1236 => (x"c2",x"87",x"f9",x"c0"),
  1237 => (x"48",x"bf",x"d8",x"eb"),
  1238 => (x"eb",x"c2",x"80",x"c1"),
  1239 => (x"eb",x"c0",x"58",x"dc"),
  1240 => (x"d8",x"eb",x"c2",x"87"),
  1241 => (x"89",x"c6",x"49",x"bf"),
  1242 => (x"59",x"dc",x"eb",x"c2"),
  1243 => (x"03",x"a9",x"b7",x"c0"),
  1244 => (x"eb",x"c2",x"87",x"da"),
  1245 => (x"78",x"c0",x"48",x"d8"),
  1246 => (x"eb",x"c2",x"87",x"d2"),
  1247 => (x"cb",x"02",x"bf",x"dc"),
  1248 => (x"d8",x"eb",x"c2",x"87"),
  1249 => (x"80",x"c6",x"48",x"bf"),
  1250 => (x"58",x"dc",x"eb",x"c2"),
  1251 => (x"f7",x"d1",x"49",x"c0"),
  1252 => (x"c0",x"49",x"73",x"87"),
  1253 => (x"f0",x"87",x"de",x"f5"),
  1254 => (x"5e",x"0e",x"87",x"dd"),
  1255 => (x"0e",x"5d",x"5c",x"5b"),
  1256 => (x"dc",x"86",x"d0",x"ff"),
  1257 => (x"a6",x"c8",x"59",x"a6"),
  1258 => (x"c4",x"78",x"c0",x"48"),
  1259 => (x"66",x"c4",x"c1",x"80"),
  1260 => (x"c1",x"80",x"c4",x"78"),
  1261 => (x"c1",x"80",x"c4",x"78"),
  1262 => (x"dc",x"eb",x"c2",x"78"),
  1263 => (x"c2",x"78",x"c1",x"48"),
  1264 => (x"48",x"bf",x"c0",x"eb"),
  1265 => (x"cb",x"05",x"a8",x"de"),
  1266 => (x"87",x"db",x"f4",x"87"),
  1267 => (x"a6",x"cc",x"49",x"70"),
  1268 => (x"87",x"f3",x"cf",x"59"),
  1269 => (x"e4",x"87",x"f7",x"e3"),
  1270 => (x"e6",x"e3",x"87",x"d9"),
  1271 => (x"c0",x"4c",x"70",x"87"),
  1272 => (x"c1",x"02",x"ac",x"fb"),
  1273 => (x"66",x"d8",x"87",x"fb"),
  1274 => (x"87",x"ed",x"c1",x"05"),
  1275 => (x"4a",x"66",x"c0",x"c1"),
  1276 => (x"7e",x"6a",x"82",x"c4"),
  1277 => (x"df",x"c1",x"1e",x"72"),
  1278 => (x"66",x"c4",x"48",x"fc"),
  1279 => (x"4a",x"a1",x"c8",x"49"),
  1280 => (x"aa",x"71",x"41",x"20"),
  1281 => (x"10",x"87",x"f9",x"05"),
  1282 => (x"c1",x"4a",x"26",x"51"),
  1283 => (x"c1",x"48",x"66",x"c0"),
  1284 => (x"6a",x"78",x"f5",x"c8"),
  1285 => (x"74",x"81",x"c7",x"49"),
  1286 => (x"66",x"c0",x"c1",x"51"),
  1287 => (x"c1",x"81",x"c8",x"49"),
  1288 => (x"66",x"c0",x"c1",x"51"),
  1289 => (x"c0",x"81",x"c9",x"49"),
  1290 => (x"66",x"c0",x"c1",x"51"),
  1291 => (x"c0",x"81",x"ca",x"49"),
  1292 => (x"d8",x"1e",x"c1",x"51"),
  1293 => (x"c8",x"49",x"6a",x"1e"),
  1294 => (x"87",x"cb",x"e3",x"81"),
  1295 => (x"c4",x"c1",x"86",x"c8"),
  1296 => (x"a8",x"c0",x"48",x"66"),
  1297 => (x"c8",x"87",x"c7",x"01"),
  1298 => (x"78",x"c1",x"48",x"a6"),
  1299 => (x"c4",x"c1",x"87",x"ce"),
  1300 => (x"88",x"c1",x"48",x"66"),
  1301 => (x"c3",x"58",x"a6",x"d0"),
  1302 => (x"87",x"d7",x"e2",x"87"),
  1303 => (x"c2",x"48",x"a6",x"d0"),
  1304 => (x"02",x"9c",x"74",x"78"),
  1305 => (x"c8",x"87",x"dc",x"cd"),
  1306 => (x"c8",x"c1",x"48",x"66"),
  1307 => (x"cd",x"03",x"a8",x"66"),
  1308 => (x"a6",x"dc",x"87",x"d1"),
  1309 => (x"e8",x"78",x"c0",x"48"),
  1310 => (x"e1",x"78",x"c0",x"80"),
  1311 => (x"4c",x"70",x"87",x"c5"),
  1312 => (x"05",x"ac",x"d0",x"c1"),
  1313 => (x"c4",x"87",x"d8",x"c2"),
  1314 => (x"e9",x"e3",x"7e",x"66"),
  1315 => (x"c8",x"49",x"70",x"87"),
  1316 => (x"ee",x"e0",x"59",x"a6"),
  1317 => (x"c0",x"4c",x"70",x"87"),
  1318 => (x"c1",x"05",x"ac",x"ec"),
  1319 => (x"66",x"c8",x"87",x"ec"),
  1320 => (x"c1",x"91",x"cb",x"49"),
  1321 => (x"c4",x"81",x"66",x"c0"),
  1322 => (x"4d",x"6a",x"4a",x"a1"),
  1323 => (x"c4",x"4a",x"a1",x"c8"),
  1324 => (x"c9",x"c1",x"52",x"66"),
  1325 => (x"ca",x"e0",x"79",x"f6"),
  1326 => (x"9c",x"4c",x"70",x"87"),
  1327 => (x"c0",x"87",x"d9",x"02"),
  1328 => (x"d3",x"02",x"ac",x"fb"),
  1329 => (x"ff",x"55",x"74",x"87"),
  1330 => (x"70",x"87",x"f8",x"df"),
  1331 => (x"c7",x"02",x"9c",x"4c"),
  1332 => (x"ac",x"fb",x"c0",x"87"),
  1333 => (x"87",x"ed",x"ff",x"05"),
  1334 => (x"c2",x"55",x"e0",x"c0"),
  1335 => (x"97",x"c0",x"55",x"c1"),
  1336 => (x"49",x"66",x"d8",x"7d"),
  1337 => (x"db",x"05",x"a9",x"6e"),
  1338 => (x"48",x"66",x"c8",x"87"),
  1339 => (x"04",x"a8",x"66",x"cc"),
  1340 => (x"66",x"c8",x"87",x"ca"),
  1341 => (x"cc",x"80",x"c1",x"48"),
  1342 => (x"87",x"c8",x"58",x"a6"),
  1343 => (x"c1",x"48",x"66",x"cc"),
  1344 => (x"58",x"a6",x"d0",x"88"),
  1345 => (x"87",x"fb",x"de",x"ff"),
  1346 => (x"d0",x"c1",x"4c",x"70"),
  1347 => (x"87",x"c8",x"05",x"ac"),
  1348 => (x"c1",x"48",x"66",x"d4"),
  1349 => (x"58",x"a6",x"d8",x"80"),
  1350 => (x"02",x"ac",x"d0",x"c1"),
  1351 => (x"c0",x"87",x"e8",x"fd"),
  1352 => (x"d8",x"48",x"a6",x"e0"),
  1353 => (x"66",x"c4",x"78",x"66"),
  1354 => (x"66",x"e0",x"c0",x"48"),
  1355 => (x"e4",x"c9",x"05",x"a8"),
  1356 => (x"a6",x"e4",x"c0",x"87"),
  1357 => (x"c4",x"78",x"c0",x"48"),
  1358 => (x"74",x"78",x"c0",x"80"),
  1359 => (x"88",x"fb",x"c0",x"48"),
  1360 => (x"02",x"6e",x"7e",x"70"),
  1361 => (x"6e",x"87",x"e7",x"c8"),
  1362 => (x"70",x"88",x"cb",x"48"),
  1363 => (x"c1",x"02",x"6e",x"7e"),
  1364 => (x"48",x"6e",x"87",x"cd"),
  1365 => (x"7e",x"70",x"88",x"c9"),
  1366 => (x"e9",x"c3",x"02",x"6e"),
  1367 => (x"c4",x"48",x"6e",x"87"),
  1368 => (x"6e",x"7e",x"70",x"88"),
  1369 => (x"6e",x"87",x"ce",x"02"),
  1370 => (x"70",x"88",x"c1",x"48"),
  1371 => (x"c3",x"02",x"6e",x"7e"),
  1372 => (x"f3",x"c7",x"87",x"d4"),
  1373 => (x"48",x"a6",x"dc",x"87"),
  1374 => (x"ff",x"78",x"f0",x"c0"),
  1375 => (x"70",x"87",x"c4",x"dd"),
  1376 => (x"ac",x"ec",x"c0",x"4c"),
  1377 => (x"87",x"c4",x"c0",x"02"),
  1378 => (x"5c",x"a6",x"e0",x"c0"),
  1379 => (x"02",x"ac",x"ec",x"c0"),
  1380 => (x"dc",x"ff",x"87",x"cd"),
  1381 => (x"4c",x"70",x"87",x"ed"),
  1382 => (x"05",x"ac",x"ec",x"c0"),
  1383 => (x"c0",x"87",x"f3",x"ff"),
  1384 => (x"c0",x"02",x"ac",x"ec"),
  1385 => (x"dc",x"ff",x"87",x"c4"),
  1386 => (x"1e",x"c0",x"87",x"d9"),
  1387 => (x"66",x"d0",x"1e",x"ca"),
  1388 => (x"c1",x"91",x"cb",x"49"),
  1389 => (x"71",x"48",x"66",x"c8"),
  1390 => (x"58",x"a6",x"cc",x"80"),
  1391 => (x"c4",x"48",x"66",x"c8"),
  1392 => (x"58",x"a6",x"d0",x"80"),
  1393 => (x"49",x"bf",x"66",x"cc"),
  1394 => (x"87",x"fb",x"dc",x"ff"),
  1395 => (x"1e",x"de",x"1e",x"c1"),
  1396 => (x"49",x"bf",x"66",x"d4"),
  1397 => (x"87",x"ef",x"dc",x"ff"),
  1398 => (x"49",x"70",x"86",x"d0"),
  1399 => (x"c0",x"89",x"09",x"c0"),
  1400 => (x"c0",x"59",x"a6",x"ec"),
  1401 => (x"c0",x"48",x"66",x"e8"),
  1402 => (x"ee",x"c0",x"06",x"a8"),
  1403 => (x"66",x"e8",x"c0",x"87"),
  1404 => (x"03",x"a8",x"dd",x"48"),
  1405 => (x"c4",x"87",x"e4",x"c0"),
  1406 => (x"c0",x"49",x"bf",x"66"),
  1407 => (x"c0",x"81",x"66",x"e8"),
  1408 => (x"e8",x"c0",x"51",x"e0"),
  1409 => (x"81",x"c1",x"49",x"66"),
  1410 => (x"81",x"bf",x"66",x"c4"),
  1411 => (x"c0",x"51",x"c1",x"c2"),
  1412 => (x"c2",x"49",x"66",x"e8"),
  1413 => (x"bf",x"66",x"c4",x"81"),
  1414 => (x"6e",x"51",x"c0",x"81"),
  1415 => (x"f5",x"c8",x"c1",x"48"),
  1416 => (x"c8",x"49",x"6e",x"78"),
  1417 => (x"51",x"66",x"d0",x"81"),
  1418 => (x"81",x"c9",x"49",x"6e"),
  1419 => (x"6e",x"51",x"66",x"d4"),
  1420 => (x"dc",x"81",x"ca",x"49"),
  1421 => (x"66",x"d0",x"51",x"66"),
  1422 => (x"d4",x"80",x"c1",x"48"),
  1423 => (x"d8",x"48",x"58",x"a6"),
  1424 => (x"c4",x"78",x"c1",x"80"),
  1425 => (x"dc",x"ff",x"87",x"e8"),
  1426 => (x"49",x"70",x"87",x"ec"),
  1427 => (x"59",x"a6",x"ec",x"c0"),
  1428 => (x"87",x"e2",x"dc",x"ff"),
  1429 => (x"e0",x"c0",x"49",x"70"),
  1430 => (x"66",x"dc",x"59",x"a6"),
  1431 => (x"a8",x"ec",x"c0",x"48"),
  1432 => (x"87",x"ca",x"c0",x"05"),
  1433 => (x"c0",x"48",x"a6",x"dc"),
  1434 => (x"c0",x"78",x"66",x"e8"),
  1435 => (x"d9",x"ff",x"87",x"c4"),
  1436 => (x"66",x"c8",x"87",x"d1"),
  1437 => (x"c1",x"91",x"cb",x"49"),
  1438 => (x"71",x"48",x"66",x"c0"),
  1439 => (x"6e",x"7e",x"70",x"80"),
  1440 => (x"6e",x"82",x"c8",x"4a"),
  1441 => (x"c0",x"81",x"ca",x"49"),
  1442 => (x"dc",x"51",x"66",x"e8"),
  1443 => (x"81",x"c1",x"49",x"66"),
  1444 => (x"89",x"66",x"e8",x"c0"),
  1445 => (x"30",x"71",x"48",x"c1"),
  1446 => (x"89",x"c1",x"49",x"70"),
  1447 => (x"c2",x"7a",x"97",x"71"),
  1448 => (x"49",x"bf",x"c8",x"ef"),
  1449 => (x"29",x"66",x"e8",x"c0"),
  1450 => (x"48",x"4a",x"6a",x"97"),
  1451 => (x"f0",x"c0",x"98",x"71"),
  1452 => (x"49",x"6e",x"58",x"a6"),
  1453 => (x"4d",x"69",x"81",x"c4"),
  1454 => (x"48",x"66",x"e0",x"c0"),
  1455 => (x"02",x"a8",x"66",x"c4"),
  1456 => (x"c4",x"87",x"c8",x"c0"),
  1457 => (x"78",x"c0",x"48",x"a6"),
  1458 => (x"c4",x"87",x"c5",x"c0"),
  1459 => (x"78",x"c1",x"48",x"a6"),
  1460 => (x"c0",x"1e",x"66",x"c4"),
  1461 => (x"49",x"75",x"1e",x"e0"),
  1462 => (x"87",x"eb",x"d8",x"ff"),
  1463 => (x"4c",x"70",x"86",x"c8"),
  1464 => (x"06",x"ac",x"b7",x"c0"),
  1465 => (x"74",x"87",x"d4",x"c1"),
  1466 => (x"49",x"e0",x"c0",x"85"),
  1467 => (x"4b",x"75",x"89",x"74"),
  1468 => (x"4a",x"c5",x"e0",x"c1"),
  1469 => (x"ef",x"e6",x"fe",x"71"),
  1470 => (x"c0",x"85",x"c2",x"87"),
  1471 => (x"c1",x"48",x"66",x"e4"),
  1472 => (x"a6",x"e8",x"c0",x"80"),
  1473 => (x"66",x"ec",x"c0",x"58"),
  1474 => (x"70",x"81",x"c1",x"49"),
  1475 => (x"c8",x"c0",x"02",x"a9"),
  1476 => (x"48",x"a6",x"c4",x"87"),
  1477 => (x"c5",x"c0",x"78",x"c0"),
  1478 => (x"48",x"a6",x"c4",x"87"),
  1479 => (x"66",x"c4",x"78",x"c1"),
  1480 => (x"49",x"a4",x"c2",x"1e"),
  1481 => (x"71",x"48",x"e0",x"c0"),
  1482 => (x"1e",x"49",x"70",x"88"),
  1483 => (x"d7",x"ff",x"49",x"75"),
  1484 => (x"86",x"c8",x"87",x"d5"),
  1485 => (x"01",x"a8",x"b7",x"c0"),
  1486 => (x"c0",x"87",x"c0",x"ff"),
  1487 => (x"c0",x"02",x"66",x"e4"),
  1488 => (x"49",x"6e",x"87",x"d1"),
  1489 => (x"e4",x"c0",x"81",x"c9"),
  1490 => (x"48",x"6e",x"51",x"66"),
  1491 => (x"78",x"c6",x"cb",x"c1"),
  1492 => (x"6e",x"87",x"cc",x"c0"),
  1493 => (x"c2",x"81",x"c9",x"49"),
  1494 => (x"c1",x"48",x"6e",x"51"),
  1495 => (x"c0",x"78",x"fa",x"cb"),
  1496 => (x"c1",x"48",x"a6",x"e8"),
  1497 => (x"87",x"c6",x"c0",x"78"),
  1498 => (x"87",x"c7",x"d6",x"ff"),
  1499 => (x"e8",x"c0",x"4c",x"70"),
  1500 => (x"f5",x"c0",x"02",x"66"),
  1501 => (x"48",x"66",x"c8",x"87"),
  1502 => (x"04",x"a8",x"66",x"cc"),
  1503 => (x"c8",x"87",x"cb",x"c0"),
  1504 => (x"80",x"c1",x"48",x"66"),
  1505 => (x"c0",x"58",x"a6",x"cc"),
  1506 => (x"66",x"cc",x"87",x"e0"),
  1507 => (x"d0",x"88",x"c1",x"48"),
  1508 => (x"d5",x"c0",x"58",x"a6"),
  1509 => (x"ac",x"c6",x"c1",x"87"),
  1510 => (x"87",x"c8",x"c0",x"05"),
  1511 => (x"c1",x"48",x"66",x"d0"),
  1512 => (x"58",x"a6",x"d4",x"80"),
  1513 => (x"87",x"cb",x"d5",x"ff"),
  1514 => (x"66",x"d4",x"4c",x"70"),
  1515 => (x"d8",x"80",x"c1",x"48"),
  1516 => (x"9c",x"74",x"58",x"a6"),
  1517 => (x"87",x"cb",x"c0",x"02"),
  1518 => (x"c1",x"48",x"66",x"c8"),
  1519 => (x"04",x"a8",x"66",x"c8"),
  1520 => (x"ff",x"87",x"ef",x"f2"),
  1521 => (x"c8",x"87",x"e3",x"d4"),
  1522 => (x"a8",x"c7",x"48",x"66"),
  1523 => (x"87",x"e5",x"c0",x"03"),
  1524 => (x"48",x"dc",x"eb",x"c2"),
  1525 => (x"66",x"c8",x"78",x"c0"),
  1526 => (x"c1",x"91",x"cb",x"49"),
  1527 => (x"c4",x"81",x"66",x"c0"),
  1528 => (x"4a",x"6a",x"4a",x"a1"),
  1529 => (x"c8",x"79",x"52",x"c0"),
  1530 => (x"80",x"c1",x"48",x"66"),
  1531 => (x"c7",x"58",x"a6",x"cc"),
  1532 => (x"db",x"ff",x"04",x"a8"),
  1533 => (x"8e",x"d0",x"ff",x"87"),
  1534 => (x"87",x"f7",x"de",x"ff"),
  1535 => (x"64",x"61",x"6f",x"4c"),
  1536 => (x"20",x"2e",x"2a",x"20"),
  1537 => (x"00",x"20",x"3a",x"00"),
  1538 => (x"71",x"1e",x"73",x"1e"),
  1539 => (x"c6",x"02",x"9b",x"4b"),
  1540 => (x"d8",x"eb",x"c2",x"87"),
  1541 => (x"c7",x"78",x"c0",x"48"),
  1542 => (x"d8",x"eb",x"c2",x"1e"),
  1543 => (x"c1",x"1e",x"49",x"bf"),
  1544 => (x"c2",x"1e",x"e4",x"e3"),
  1545 => (x"49",x"bf",x"c0",x"eb"),
  1546 => (x"cc",x"87",x"ef",x"ed"),
  1547 => (x"c0",x"eb",x"c2",x"86"),
  1548 => (x"e9",x"e9",x"49",x"bf"),
  1549 => (x"02",x"9b",x"73",x"87"),
  1550 => (x"e3",x"c1",x"87",x"c8"),
  1551 => (x"e4",x"c0",x"49",x"e4"),
  1552 => (x"dd",x"ff",x"87",x"c5"),
  1553 => (x"c7",x"1e",x"87",x"f1"),
  1554 => (x"49",x"c1",x"87",x"d4"),
  1555 => (x"fe",x"87",x"f9",x"fe"),
  1556 => (x"70",x"87",x"fd",x"e9"),
  1557 => (x"87",x"cd",x"02",x"98"),
  1558 => (x"87",x"f8",x"f2",x"fe"),
  1559 => (x"c4",x"02",x"98",x"70"),
  1560 => (x"c2",x"4a",x"c1",x"87"),
  1561 => (x"72",x"4a",x"c0",x"87"),
  1562 => (x"87",x"ce",x"05",x"9a"),
  1563 => (x"e2",x"c1",x"1e",x"c0"),
  1564 => (x"ef",x"c0",x"49",x"d7"),
  1565 => (x"86",x"c4",x"87",x"e0"),
  1566 => (x"1e",x"c0",x"87",x"fe"),
  1567 => (x"49",x"e2",x"e2",x"c1"),
  1568 => (x"87",x"d2",x"ef",x"c0"),
  1569 => (x"f9",x"c0",x"1e",x"c0"),
  1570 => (x"49",x"70",x"87",x"c0"),
  1571 => (x"87",x"c6",x"ef",x"c0"),
  1572 => (x"f8",x"87",x"ca",x"c3"),
  1573 => (x"53",x"4f",x"26",x"8e"),
  1574 => (x"61",x"66",x"20",x"44"),
  1575 => (x"64",x"65",x"6c",x"69"),
  1576 => (x"6f",x"42",x"00",x"2e"),
  1577 => (x"6e",x"69",x"74",x"6f"),
  1578 => (x"2e",x"2e",x"2e",x"67"),
  1579 => (x"e6",x"c0",x"1e",x"00"),
  1580 => (x"f2",x"c0",x"87",x"f1"),
  1581 => (x"87",x"f6",x"87",x"d6"),
  1582 => (x"c2",x"1e",x"4f",x"26"),
  1583 => (x"c0",x"48",x"d8",x"eb"),
  1584 => (x"c0",x"eb",x"c2",x"78"),
  1585 => (x"fd",x"78",x"c0",x"48"),
  1586 => (x"87",x"e1",x"87",x"fc"),
  1587 => (x"4f",x"26",x"48",x"c0"),
  1588 => (x"00",x"01",x"00",x"00"),
  1589 => (x"20",x"80",x"00",x"00"),
  1590 => (x"74",x"69",x"78",x"45"),
  1591 => (x"42",x"20",x"80",x"00"),
  1592 => (x"00",x"6b",x"63",x"61"),
  1593 => (x"00",x"00",x"12",x"76"),
  1594 => (x"00",x"00",x"2a",x"ec"),
  1595 => (x"76",x"00",x"00",x"00"),
  1596 => (x"0a",x"00",x"00",x"12"),
  1597 => (x"00",x"00",x"00",x"2b"),
  1598 => (x"12",x"76",x"00",x"00"),
  1599 => (x"2b",x"28",x"00",x"00"),
  1600 => (x"00",x"00",x"00",x"00"),
  1601 => (x"00",x"12",x"76",x"00"),
  1602 => (x"00",x"2b",x"46",x"00"),
  1603 => (x"00",x"00",x"00",x"00"),
  1604 => (x"00",x"00",x"12",x"76"),
  1605 => (x"00",x"00",x"2b",x"64"),
  1606 => (x"76",x"00",x"00",x"00"),
  1607 => (x"82",x"00",x"00",x"12"),
  1608 => (x"00",x"00",x"00",x"2b"),
  1609 => (x"12",x"76",x"00",x"00"),
  1610 => (x"2b",x"a0",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"12",x"76",x"00"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"13",x"0b"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"1e",x"00",x"00",x"00"),
  1618 => (x"c0",x"48",x"f0",x"fe"),
  1619 => (x"79",x"09",x"cd",x"78"),
  1620 => (x"1e",x"4f",x"26",x"09"),
  1621 => (x"bf",x"f0",x"fe",x"1e"),
  1622 => (x"26",x"26",x"48",x"7e"),
  1623 => (x"f0",x"fe",x"1e",x"4f"),
  1624 => (x"26",x"78",x"c1",x"48"),
  1625 => (x"f0",x"fe",x"1e",x"4f"),
  1626 => (x"26",x"78",x"c0",x"48"),
  1627 => (x"4a",x"71",x"1e",x"4f"),
  1628 => (x"26",x"52",x"52",x"c0"),
  1629 => (x"5b",x"5e",x"0e",x"4f"),
  1630 => (x"f4",x"0e",x"5d",x"5c"),
  1631 => (x"97",x"4d",x"71",x"86"),
  1632 => (x"a5",x"c1",x"7e",x"6d"),
  1633 => (x"48",x"6c",x"97",x"4c"),
  1634 => (x"6e",x"58",x"a6",x"c8"),
  1635 => (x"a8",x"66",x"c4",x"48"),
  1636 => (x"ff",x"87",x"c5",x"05"),
  1637 => (x"87",x"e6",x"c0",x"48"),
  1638 => (x"c2",x"87",x"ca",x"ff"),
  1639 => (x"6c",x"97",x"49",x"a5"),
  1640 => (x"4b",x"a3",x"71",x"4b"),
  1641 => (x"97",x"4b",x"6b",x"97"),
  1642 => (x"48",x"6e",x"7e",x"6c"),
  1643 => (x"a6",x"c8",x"80",x"c1"),
  1644 => (x"cc",x"98",x"c7",x"58"),
  1645 => (x"97",x"70",x"58",x"a6"),
  1646 => (x"87",x"e1",x"fe",x"7c"),
  1647 => (x"8e",x"f4",x"48",x"73"),
  1648 => (x"4c",x"26",x"4d",x"26"),
  1649 => (x"4f",x"26",x"4b",x"26"),
  1650 => (x"5c",x"5b",x"5e",x"0e"),
  1651 => (x"71",x"86",x"f4",x"0e"),
  1652 => (x"4a",x"66",x"d8",x"4c"),
  1653 => (x"c2",x"9a",x"ff",x"c3"),
  1654 => (x"6c",x"97",x"4b",x"a4"),
  1655 => (x"49",x"a1",x"73",x"49"),
  1656 => (x"6c",x"97",x"51",x"72"),
  1657 => (x"c1",x"48",x"6e",x"7e"),
  1658 => (x"58",x"a6",x"c8",x"80"),
  1659 => (x"a6",x"cc",x"98",x"c7"),
  1660 => (x"f4",x"54",x"70",x"58"),
  1661 => (x"87",x"ca",x"ff",x"8e"),
  1662 => (x"e8",x"fd",x"1e",x"1e"),
  1663 => (x"4a",x"bf",x"e0",x"87"),
  1664 => (x"c0",x"e0",x"c0",x"49"),
  1665 => (x"87",x"cb",x"02",x"99"),
  1666 => (x"ee",x"c2",x"1e",x"72"),
  1667 => (x"f7",x"fe",x"49",x"fe"),
  1668 => (x"fc",x"86",x"c4",x"87"),
  1669 => (x"7e",x"70",x"87",x"fd"),
  1670 => (x"26",x"87",x"c2",x"fd"),
  1671 => (x"c2",x"1e",x"4f",x"26"),
  1672 => (x"fd",x"49",x"fe",x"ee"),
  1673 => (x"e7",x"c1",x"87",x"c7"),
  1674 => (x"da",x"fc",x"49",x"f8"),
  1675 => (x"87",x"f7",x"c3",x"87"),
  1676 => (x"5e",x"0e",x"4f",x"26"),
  1677 => (x"0e",x"5d",x"5c",x"5b"),
  1678 => (x"ee",x"c2",x"4d",x"71"),
  1679 => (x"f4",x"fc",x"49",x"fe"),
  1680 => (x"c0",x"4b",x"70",x"87"),
  1681 => (x"c3",x"04",x"ab",x"b7"),
  1682 => (x"f0",x"c3",x"87",x"c2"),
  1683 => (x"87",x"c9",x"05",x"ab"),
  1684 => (x"48",x"d6",x"ec",x"c1"),
  1685 => (x"e3",x"c2",x"78",x"c1"),
  1686 => (x"ab",x"e0",x"c3",x"87"),
  1687 => (x"c1",x"87",x"c9",x"05"),
  1688 => (x"c1",x"48",x"da",x"ec"),
  1689 => (x"87",x"d4",x"c2",x"78"),
  1690 => (x"bf",x"da",x"ec",x"c1"),
  1691 => (x"c2",x"87",x"c6",x"02"),
  1692 => (x"c2",x"4c",x"a3",x"c0"),
  1693 => (x"c1",x"4c",x"73",x"87"),
  1694 => (x"02",x"bf",x"d6",x"ec"),
  1695 => (x"74",x"87",x"e0",x"c0"),
  1696 => (x"29",x"b7",x"c4",x"49"),
  1697 => (x"f6",x"ed",x"c1",x"91"),
  1698 => (x"cf",x"4a",x"74",x"81"),
  1699 => (x"c1",x"92",x"c2",x"9a"),
  1700 => (x"70",x"30",x"72",x"48"),
  1701 => (x"72",x"ba",x"ff",x"4a"),
  1702 => (x"70",x"98",x"69",x"48"),
  1703 => (x"74",x"87",x"db",x"79"),
  1704 => (x"29",x"b7",x"c4",x"49"),
  1705 => (x"f6",x"ed",x"c1",x"91"),
  1706 => (x"cf",x"4a",x"74",x"81"),
  1707 => (x"c3",x"92",x"c2",x"9a"),
  1708 => (x"70",x"30",x"72",x"48"),
  1709 => (x"b0",x"69",x"48",x"4a"),
  1710 => (x"9d",x"75",x"79",x"70"),
  1711 => (x"87",x"f0",x"c0",x"05"),
  1712 => (x"c8",x"48",x"d0",x"ff"),
  1713 => (x"d4",x"ff",x"78",x"e1"),
  1714 => (x"c1",x"78",x"c5",x"48"),
  1715 => (x"02",x"bf",x"da",x"ec"),
  1716 => (x"e0",x"c3",x"87",x"c3"),
  1717 => (x"d6",x"ec",x"c1",x"78"),
  1718 => (x"87",x"c6",x"02",x"bf"),
  1719 => (x"c3",x"48",x"d4",x"ff"),
  1720 => (x"d4",x"ff",x"78",x"f0"),
  1721 => (x"ff",x"78",x"73",x"48"),
  1722 => (x"e1",x"c8",x"48",x"d0"),
  1723 => (x"78",x"e0",x"c0",x"78"),
  1724 => (x"48",x"da",x"ec",x"c1"),
  1725 => (x"ec",x"c1",x"78",x"c0"),
  1726 => (x"78",x"c0",x"48",x"d6"),
  1727 => (x"49",x"fe",x"ee",x"c2"),
  1728 => (x"70",x"87",x"f2",x"f9"),
  1729 => (x"ab",x"b7",x"c0",x"4b"),
  1730 => (x"87",x"fe",x"fc",x"03"),
  1731 => (x"4d",x"26",x"48",x"c0"),
  1732 => (x"4b",x"26",x"4c",x"26"),
  1733 => (x"00",x"00",x"4f",x"26"),
  1734 => (x"00",x"00",x"00",x"00"),
  1735 => (x"71",x"1e",x"00",x"00"),
  1736 => (x"cd",x"fc",x"49",x"4a"),
  1737 => (x"1e",x"4f",x"26",x"87"),
  1738 => (x"49",x"72",x"4a",x"c0"),
  1739 => (x"ed",x"c1",x"91",x"c4"),
  1740 => (x"79",x"c0",x"81",x"f6"),
  1741 => (x"b7",x"d0",x"82",x"c1"),
  1742 => (x"87",x"ee",x"04",x"aa"),
  1743 => (x"5e",x"0e",x"4f",x"26"),
  1744 => (x"0e",x"5d",x"5c",x"5b"),
  1745 => (x"dc",x"f8",x"4d",x"71"),
  1746 => (x"c4",x"4a",x"75",x"87"),
  1747 => (x"c1",x"92",x"2a",x"b7"),
  1748 => (x"75",x"82",x"f6",x"ed"),
  1749 => (x"c2",x"9c",x"cf",x"4c"),
  1750 => (x"4b",x"49",x"6a",x"94"),
  1751 => (x"9b",x"c3",x"2b",x"74"),
  1752 => (x"30",x"74",x"48",x"c2"),
  1753 => (x"bc",x"ff",x"4c",x"70"),
  1754 => (x"98",x"71",x"48",x"74"),
  1755 => (x"ec",x"f7",x"7a",x"70"),
  1756 => (x"fe",x"48",x"73",x"87"),
  1757 => (x"00",x"00",x"87",x"d8"),
  1758 => (x"40",x"40",x"00",x"00"),
  1759 => (x"40",x"40",x"40",x"40"),
  1760 => (x"40",x"40",x"40",x"40"),
  1761 => (x"40",x"40",x"40",x"40"),
  1762 => (x"40",x"40",x"40",x"40"),
  1763 => (x"40",x"40",x"40",x"40"),
  1764 => (x"40",x"40",x"40",x"40"),
  1765 => (x"40",x"40",x"40",x"40"),
  1766 => (x"40",x"40",x"40",x"40"),
  1767 => (x"40",x"40",x"40",x"40"),
  1768 => (x"40",x"40",x"40",x"40"),
  1769 => (x"40",x"40",x"40",x"40"),
  1770 => (x"40",x"40",x"40",x"40"),
  1771 => (x"40",x"40",x"40",x"40"),
  1772 => (x"40",x"40",x"40",x"40"),
  1773 => (x"ff",x"1e",x"40",x"40"),
  1774 => (x"e1",x"c8",x"48",x"d0"),
  1775 => (x"ff",x"48",x"71",x"78"),
  1776 => (x"26",x"78",x"08",x"d4"),
  1777 => (x"d0",x"ff",x"1e",x"4f"),
  1778 => (x"78",x"e1",x"c8",x"48"),
  1779 => (x"d4",x"ff",x"48",x"71"),
  1780 => (x"66",x"c4",x"78",x"08"),
  1781 => (x"08",x"d4",x"ff",x"48"),
  1782 => (x"1e",x"4f",x"26",x"78"),
  1783 => (x"66",x"c4",x"4a",x"71"),
  1784 => (x"49",x"72",x"1e",x"49"),
  1785 => (x"ff",x"87",x"de",x"ff"),
  1786 => (x"e0",x"c0",x"48",x"d0"),
  1787 => (x"4f",x"26",x"26",x"78"),
  1788 => (x"71",x"1e",x"73",x"1e"),
  1789 => (x"49",x"66",x"c8",x"4b"),
  1790 => (x"c1",x"4a",x"73",x"1e"),
  1791 => (x"ff",x"49",x"a2",x"e0"),
  1792 => (x"c4",x"26",x"87",x"d9"),
  1793 => (x"26",x"4d",x"26",x"87"),
  1794 => (x"26",x"4b",x"26",x"4c"),
  1795 => (x"1e",x"73",x"1e",x"4f"),
  1796 => (x"c2",x"4b",x"4a",x"71"),
  1797 => (x"c8",x"03",x"ab",x"b7"),
  1798 => (x"4a",x"49",x"a3",x"87"),
  1799 => (x"c7",x"9a",x"ff",x"c3"),
  1800 => (x"49",x"a3",x"ce",x"87"),
  1801 => (x"9a",x"ff",x"c3",x"4a"),
  1802 => (x"1e",x"49",x"66",x"c8"),
  1803 => (x"ea",x"fe",x"49",x"72"),
  1804 => (x"d4",x"ff",x"26",x"87"),
  1805 => (x"d4",x"ff",x"1e",x"87"),
  1806 => (x"7a",x"ff",x"c3",x"4a"),
  1807 => (x"c0",x"48",x"d0",x"ff"),
  1808 => (x"7a",x"de",x"78",x"e1"),
  1809 => (x"bf",x"c8",x"ef",x"c2"),
  1810 => (x"c8",x"48",x"49",x"7a"),
  1811 => (x"71",x"7a",x"70",x"28"),
  1812 => (x"70",x"28",x"d0",x"48"),
  1813 => (x"d8",x"48",x"71",x"7a"),
  1814 => (x"ff",x"7a",x"70",x"28"),
  1815 => (x"e0",x"c0",x"48",x"d0"),
  1816 => (x"0e",x"4f",x"26",x"78"),
  1817 => (x"5d",x"5c",x"5b",x"5e"),
  1818 => (x"c2",x"4c",x"71",x"0e"),
  1819 => (x"4d",x"bf",x"c8",x"ef"),
  1820 => (x"71",x"29",x"74",x"49"),
  1821 => (x"9b",x"66",x"d0",x"4b"),
  1822 => (x"66",x"d4",x"83",x"c1"),
  1823 => (x"c2",x"04",x"ab",x"b7"),
  1824 => (x"d0",x"4b",x"c0",x"87"),
  1825 => (x"31",x"74",x"49",x"66"),
  1826 => (x"99",x"75",x"b9",x"ff"),
  1827 => (x"32",x"74",x"4a",x"73"),
  1828 => (x"b0",x"71",x"48",x"72"),
  1829 => (x"58",x"cc",x"ef",x"c2"),
  1830 => (x"26",x"87",x"da",x"fe"),
  1831 => (x"26",x"4c",x"26",x"4d"),
  1832 => (x"1e",x"4f",x"26",x"4b"),
  1833 => (x"c8",x"48",x"d0",x"ff"),
  1834 => (x"48",x"71",x"78",x"c9"),
  1835 => (x"78",x"08",x"d4",x"ff"),
  1836 => (x"71",x"1e",x"4f",x"26"),
  1837 => (x"87",x"eb",x"49",x"4a"),
  1838 => (x"c8",x"48",x"d0",x"ff"),
  1839 => (x"1e",x"4f",x"26",x"78"),
  1840 => (x"4b",x"71",x"1e",x"73"),
  1841 => (x"bf",x"d8",x"ef",x"c2"),
  1842 => (x"c2",x"87",x"c3",x"02"),
  1843 => (x"d0",x"ff",x"87",x"eb"),
  1844 => (x"78",x"c9",x"c8",x"48"),
  1845 => (x"e0",x"c0",x"49",x"73"),
  1846 => (x"48",x"d4",x"ff",x"b1"),
  1847 => (x"ef",x"c2",x"78",x"71"),
  1848 => (x"78",x"c0",x"48",x"cc"),
  1849 => (x"c5",x"02",x"66",x"c8"),
  1850 => (x"49",x"ff",x"c3",x"87"),
  1851 => (x"49",x"c0",x"87",x"c2"),
  1852 => (x"59",x"d4",x"ef",x"c2"),
  1853 => (x"c6",x"02",x"66",x"cc"),
  1854 => (x"d5",x"d5",x"c5",x"87"),
  1855 => (x"cf",x"87",x"c4",x"4a"),
  1856 => (x"c2",x"4a",x"ff",x"ff"),
  1857 => (x"c2",x"5a",x"d8",x"ef"),
  1858 => (x"c1",x"48",x"d8",x"ef"),
  1859 => (x"26",x"87",x"c4",x"78"),
  1860 => (x"26",x"4c",x"26",x"4d"),
  1861 => (x"0e",x"4f",x"26",x"4b"),
  1862 => (x"5d",x"5c",x"5b",x"5e"),
  1863 => (x"c2",x"4a",x"71",x"0e"),
  1864 => (x"4c",x"bf",x"d4",x"ef"),
  1865 => (x"cb",x"02",x"9a",x"72"),
  1866 => (x"91",x"c8",x"49",x"87"),
  1867 => (x"4b",x"f5",x"f2",x"c1"),
  1868 => (x"87",x"c4",x"83",x"71"),
  1869 => (x"4b",x"f5",x"f6",x"c1"),
  1870 => (x"49",x"13",x"4d",x"c0"),
  1871 => (x"ef",x"c2",x"99",x"74"),
  1872 => (x"ff",x"b9",x"bf",x"d0"),
  1873 => (x"78",x"71",x"48",x"d4"),
  1874 => (x"85",x"2c",x"b7",x"c1"),
  1875 => (x"04",x"ad",x"b7",x"c8"),
  1876 => (x"ef",x"c2",x"87",x"e8"),
  1877 => (x"c8",x"48",x"bf",x"cc"),
  1878 => (x"d0",x"ef",x"c2",x"80"),
  1879 => (x"87",x"ef",x"fe",x"58"),
  1880 => (x"71",x"1e",x"73",x"1e"),
  1881 => (x"9a",x"4a",x"13",x"4b"),
  1882 => (x"72",x"87",x"cb",x"02"),
  1883 => (x"87",x"e7",x"fe",x"49"),
  1884 => (x"05",x"9a",x"4a",x"13"),
  1885 => (x"da",x"fe",x"87",x"f5"),
  1886 => (x"ef",x"c2",x"1e",x"87"),
  1887 => (x"c2",x"49",x"bf",x"cc"),
  1888 => (x"c1",x"48",x"cc",x"ef"),
  1889 => (x"c0",x"c4",x"78",x"a1"),
  1890 => (x"db",x"03",x"a9",x"b7"),
  1891 => (x"48",x"d4",x"ff",x"87"),
  1892 => (x"bf",x"d0",x"ef",x"c2"),
  1893 => (x"cc",x"ef",x"c2",x"78"),
  1894 => (x"ef",x"c2",x"49",x"bf"),
  1895 => (x"a1",x"c1",x"48",x"cc"),
  1896 => (x"b7",x"c0",x"c4",x"78"),
  1897 => (x"87",x"e5",x"04",x"a9"),
  1898 => (x"c8",x"48",x"d0",x"ff"),
  1899 => (x"d8",x"ef",x"c2",x"78"),
  1900 => (x"26",x"78",x"c0",x"48"),
  1901 => (x"00",x"00",x"00",x"4f"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"00",x"00",x"00",x"00"),
  1904 => (x"00",x"00",x"5f",x"5f"),
  1905 => (x"03",x"03",x"00",x"00"),
  1906 => (x"00",x"03",x"03",x"00"),
  1907 => (x"7f",x"7f",x"14",x"00"),
  1908 => (x"14",x"7f",x"7f",x"14"),
  1909 => (x"2e",x"24",x"00",x"00"),
  1910 => (x"12",x"3a",x"6b",x"6b"),
  1911 => (x"36",x"6a",x"4c",x"00"),
  1912 => (x"32",x"56",x"6c",x"18"),
  1913 => (x"4f",x"7e",x"30",x"00"),
  1914 => (x"68",x"3a",x"77",x"59"),
  1915 => (x"04",x"00",x"00",x"40"),
  1916 => (x"00",x"00",x"03",x"07"),
  1917 => (x"1c",x"00",x"00",x"00"),
  1918 => (x"00",x"41",x"63",x"3e"),
  1919 => (x"41",x"00",x"00",x"00"),
  1920 => (x"00",x"1c",x"3e",x"63"),
  1921 => (x"3e",x"2a",x"08",x"00"),
  1922 => (x"2a",x"3e",x"1c",x"1c"),
  1923 => (x"08",x"08",x"00",x"08"),
  1924 => (x"08",x"08",x"3e",x"3e"),
  1925 => (x"80",x"00",x"00",x"00"),
  1926 => (x"00",x"00",x"60",x"e0"),
  1927 => (x"08",x"08",x"00",x"00"),
  1928 => (x"08",x"08",x"08",x"08"),
  1929 => (x"00",x"00",x"00",x"00"),
  1930 => (x"00",x"00",x"60",x"60"),
  1931 => (x"30",x"60",x"40",x"00"),
  1932 => (x"03",x"06",x"0c",x"18"),
  1933 => (x"7f",x"3e",x"00",x"01"),
  1934 => (x"3e",x"7f",x"4d",x"59"),
  1935 => (x"06",x"04",x"00",x"00"),
  1936 => (x"00",x"00",x"7f",x"7f"),
  1937 => (x"63",x"42",x"00",x"00"),
  1938 => (x"46",x"4f",x"59",x"71"),
  1939 => (x"63",x"22",x"00",x"00"),
  1940 => (x"36",x"7f",x"49",x"49"),
  1941 => (x"16",x"1c",x"18",x"00"),
  1942 => (x"10",x"7f",x"7f",x"13"),
  1943 => (x"67",x"27",x"00",x"00"),
  1944 => (x"39",x"7d",x"45",x"45"),
  1945 => (x"7e",x"3c",x"00",x"00"),
  1946 => (x"30",x"79",x"49",x"4b"),
  1947 => (x"01",x"01",x"00",x"00"),
  1948 => (x"07",x"0f",x"79",x"71"),
  1949 => (x"7f",x"36",x"00",x"00"),
  1950 => (x"36",x"7f",x"49",x"49"),
  1951 => (x"4f",x"06",x"00",x"00"),
  1952 => (x"1e",x"3f",x"69",x"49"),
  1953 => (x"00",x"00",x"00",x"00"),
  1954 => (x"00",x"00",x"66",x"66"),
  1955 => (x"80",x"00",x"00",x"00"),
  1956 => (x"00",x"00",x"66",x"e6"),
  1957 => (x"08",x"08",x"00",x"00"),
  1958 => (x"22",x"22",x"14",x"14"),
  1959 => (x"14",x"14",x"00",x"00"),
  1960 => (x"14",x"14",x"14",x"14"),
  1961 => (x"22",x"22",x"00",x"00"),
  1962 => (x"08",x"08",x"14",x"14"),
  1963 => (x"03",x"02",x"00",x"00"),
  1964 => (x"06",x"0f",x"59",x"51"),
  1965 => (x"41",x"7f",x"3e",x"00"),
  1966 => (x"1e",x"1f",x"55",x"5d"),
  1967 => (x"7f",x"7e",x"00",x"00"),
  1968 => (x"7e",x"7f",x"09",x"09"),
  1969 => (x"7f",x"7f",x"00",x"00"),
  1970 => (x"36",x"7f",x"49",x"49"),
  1971 => (x"3e",x"1c",x"00",x"00"),
  1972 => (x"41",x"41",x"41",x"63"),
  1973 => (x"7f",x"7f",x"00",x"00"),
  1974 => (x"1c",x"3e",x"63",x"41"),
  1975 => (x"7f",x"7f",x"00",x"00"),
  1976 => (x"41",x"41",x"49",x"49"),
  1977 => (x"7f",x"7f",x"00",x"00"),
  1978 => (x"01",x"01",x"09",x"09"),
  1979 => (x"7f",x"3e",x"00",x"00"),
  1980 => (x"7a",x"7b",x"49",x"41"),
  1981 => (x"7f",x"7f",x"00",x"00"),
  1982 => (x"7f",x"7f",x"08",x"08"),
  1983 => (x"41",x"00",x"00",x"00"),
  1984 => (x"00",x"41",x"7f",x"7f"),
  1985 => (x"60",x"20",x"00",x"00"),
  1986 => (x"3f",x"7f",x"40",x"40"),
  1987 => (x"08",x"7f",x"7f",x"00"),
  1988 => (x"41",x"63",x"36",x"1c"),
  1989 => (x"7f",x"7f",x"00",x"00"),
  1990 => (x"40",x"40",x"40",x"40"),
  1991 => (x"06",x"7f",x"7f",x"00"),
  1992 => (x"7f",x"7f",x"06",x"0c"),
  1993 => (x"06",x"7f",x"7f",x"00"),
  1994 => (x"7f",x"7f",x"18",x"0c"),
  1995 => (x"7f",x"3e",x"00",x"00"),
  1996 => (x"3e",x"7f",x"41",x"41"),
  1997 => (x"7f",x"7f",x"00",x"00"),
  1998 => (x"06",x"0f",x"09",x"09"),
  1999 => (x"41",x"7f",x"3e",x"00"),
  2000 => (x"40",x"7e",x"7f",x"61"),
  2001 => (x"7f",x"7f",x"00",x"00"),
  2002 => (x"66",x"7f",x"19",x"09"),
  2003 => (x"6f",x"26",x"00",x"00"),
  2004 => (x"32",x"7b",x"59",x"4d"),
  2005 => (x"01",x"01",x"00",x"00"),
  2006 => (x"01",x"01",x"7f",x"7f"),
  2007 => (x"7f",x"3f",x"00",x"00"),
  2008 => (x"3f",x"7f",x"40",x"40"),
  2009 => (x"3f",x"0f",x"00",x"00"),
  2010 => (x"0f",x"3f",x"70",x"70"),
  2011 => (x"30",x"7f",x"7f",x"00"),
  2012 => (x"7f",x"7f",x"30",x"18"),
  2013 => (x"36",x"63",x"41",x"00"),
  2014 => (x"63",x"36",x"1c",x"1c"),
  2015 => (x"06",x"03",x"01",x"41"),
  2016 => (x"03",x"06",x"7c",x"7c"),
  2017 => (x"59",x"71",x"61",x"01"),
  2018 => (x"41",x"43",x"47",x"4d"),
  2019 => (x"7f",x"00",x"00",x"00"),
  2020 => (x"00",x"41",x"41",x"7f"),
  2021 => (x"06",x"03",x"01",x"00"),
  2022 => (x"60",x"30",x"18",x"0c"),
  2023 => (x"41",x"00",x"00",x"40"),
  2024 => (x"00",x"7f",x"7f",x"41"),
  2025 => (x"06",x"0c",x"08",x"00"),
  2026 => (x"08",x"0c",x"06",x"03"),
  2027 => (x"80",x"80",x"80",x"00"),
  2028 => (x"80",x"80",x"80",x"80"),
  2029 => (x"00",x"00",x"00",x"00"),
  2030 => (x"00",x"04",x"07",x"03"),
  2031 => (x"74",x"20",x"00",x"00"),
  2032 => (x"78",x"7c",x"54",x"54"),
  2033 => (x"7f",x"7f",x"00",x"00"),
  2034 => (x"38",x"7c",x"44",x"44"),
  2035 => (x"7c",x"38",x"00",x"00"),
  2036 => (x"00",x"44",x"44",x"44"),
  2037 => (x"7c",x"38",x"00",x"00"),
  2038 => (x"7f",x"7f",x"44",x"44"),
  2039 => (x"7c",x"38",x"00",x"00"),
  2040 => (x"18",x"5c",x"54",x"54"),
  2041 => (x"7e",x"04",x"00",x"00"),
  2042 => (x"00",x"05",x"05",x"7f"),
  2043 => (x"bc",x"18",x"00",x"00"),
  2044 => (x"7c",x"fc",x"a4",x"a4"),
  2045 => (x"7f",x"7f",x"00",x"00"),
  2046 => (x"78",x"7c",x"04",x"04"),
  2047 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

